<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-161.358,42.6019,370.877,-236.611</PageViewport>
<gate>
<ID>1</ID>
<type>DA_FROM</type>
<position>-9.5,-48.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>2</ID>
<type>DE_TO</type>
<position>-4,19</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>3</ID>
<type>DA_FROM</type>
<position>-8,-44.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>-9,19</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_INVERTER</type>
<position>-1.5,-44.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-9,15.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_AND2</type>
<position>7.5,-46.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>DE_TO</type>
<position>-4,15.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>9</ID>
<type>GA_LED</type>
<position>13.5,-43.5</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>DA_FROM</type>
<position>-9.5,-17.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>11</ID>
<type>DA_FROM</type>
<position>-8,-54</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>-8,-13.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>13</ID>
<type>DA_FROM</type>
<position>-9.5,-58</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_INVERTER</type>
<position>-0.5,-54</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND2</type>
<position>7.5,-56</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>13.5,-59.5</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>DA_FROM</type>
<position>-8,-40.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_INVERTER</type>
<position>-1.5,-13.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>19</ID>
<type>AI_XOR2</type>
<position>23.5,-45.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND2</type>
<position>7.5,-15.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>27.5,-41</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>13.5,-12.5</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>DA_FROM</type>
<position>-8,-62</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>4,19</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AI_XOR2</type>
<position>23,-59</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>-9,12</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>27,-62</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>DE_TO</type>
<position>9,19</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>36.5,-44</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>DE_TO</type>
<position>-4,12</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>41.5,-38.5</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>DA_FROM</type>
<position>-8,-23</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_FULLADDER_1BIT</type>
<position>37.5,-55.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_B_0</ID>32 </input>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>-9.5,-27</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>37.5,-63</position>
<input>
<ID>N_in3</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_INVERTER</type>
<position>-0.5,-23</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>37</ID>
<type>DA_FROM</type>
<position>-10,-51.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>7.5,-25</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_INVERTER</type>
<position>44.5,-48.5</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>13.5,-28.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>52,-41</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>4,12</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_AND2</type>
<position>52,-56</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>4,15.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_OR2</type>
<position>61.5,-48</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>9,15.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>56,-39</position>
<input>
<ID>N_in2</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>9,12</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>49</ID>
<type>GA_LED</type>
<position>56,-61</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>DA_FROM</type>
<position>-8,-9.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>51</ID>
<type>DA_FROM</type>
<position>-8,-36.5</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>52</ID>
<type>AI_XOR2</type>
<position>23.5,-14.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AI_XOR2</type>
<position>72.5,-48</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>65.5,-52.5</position>
<input>
<ID>N_in3</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>GA_LED</type>
<position>78.5,-48</position>
<input>
<ID>N_in0</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>27.5,-10</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AE_OR2</type>
<position>78.5,-54.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>-8,-31</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>76,-59</position>
<input>
<ID>N_in3</ID>54 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AI_XOR2</type>
<position>23,-28</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_INVERTER</type>
<position>88,-54.5</position>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>92,-54.5</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>-10,-78.5</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>27,-31</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>-8.5,-74.5</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_AND2</type>
<position>36.5,-13</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_INVERTER</type>
<position>-2,-74.5</position>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>68</ID>
<type>GA_LED</type>
<position>41.5,-7.5</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>7,-76.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_FULLADDER_1BIT</type>
<position>37.5,-24.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_B_0</ID>20 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>71</ID>
<type>GA_LED</type>
<position>13,-73.5</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>GA_LED</type>
<position>37.5,-32</position>
<input>
<ID>N_in3</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>DA_FROM</type>
<position>-8.5,-84</position>
<input>
<ID>IN_0</ID>58 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>74</ID>
<type>DE_TO</type>
<position>22.5,15.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>75</ID>
<type>DA_FROM</type>
<position>-10,-88</position>
<input>
<ID>IN_0</ID>60 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>17,15.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_INVERTER</type>
<position>-1,-84</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>-10,-20.5</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>7,-86</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_INVERTER</type>
<position>44.5,-17.5</position>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>13,-89.5</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>52,-10</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>-8.5,-70.5</position>
<input>
<ID>IN_0</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_AND2</type>
<position>52,-25</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AI_XOR2</type>
<position>23,-75.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_OR2</type>
<position>61.5,-17</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>GA_LED</type>
<position>27,-71</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>56,-8</position>
<input>
<ID>N_in2</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>DA_FROM</type>
<position>-8.5,-92</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>56,-30</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AI_XOR2</type>
<position>22.5,-89</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>DE_TO</type>
<position>35,15.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>93</ID>
<type>GA_LED</type>
<position>26.5,-92</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>29,15.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_AND2</type>
<position>36,-74</position>
<input>
<ID>IN_0</ID>64 </input>
<input>
<ID>IN_1</ID>66 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>41,-68.5</position>
<input>
<ID>N_in0</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_FULLADDER_1BIT</type>
<position>37,-85.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_B_0</ID>64 </input>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>98</ID>
<type>GA_LED</type>
<position>37,-93</position>
<input>
<ID>N_in3</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>DA_FROM</type>
<position>-10.5,-81.5</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>100</ID>
<type>DA_FROM</type>
<position>-8,-5.5</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_INVERTER</type>
<position>44,-78.5</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>102</ID>
<type>AI_XOR2</type>
<position>72.5,-17</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND2</type>
<position>51.5,-71</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>GA_LED</type>
<position>65.5,-21.5</position>
<input>
<ID>N_in3</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND2</type>
<position>51.5,-86</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AE_OR2</type>
<position>61,-78</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>68 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>GA_LED</type>
<position>55.5,-69</position>
<input>
<ID>N_in2</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>GA_LED</type>
<position>55.5,-91</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>DA_FROM</type>
<position>-8.5,-66.5</position>
<input>
<ID>IN_0</ID>74 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>110</ID>
<type>GA_LED</type>
<position>78.5,-17</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AI_XOR2</type>
<position>72,-78</position>
<input>
<ID>IN_0</ID>74 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AE_OR2</type>
<position>78.5,-23.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>GA_LED</type>
<position>65,-82.5</position>
<input>
<ID>N_in3</ID>69 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>GA_LED</type>
<position>76,-28</position>
<input>
<ID>N_in3</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>78,-78</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_INVERTER</type>
<position>88,-23.5</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_OR2</type>
<position>78,-84.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>77 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>GA_LED</type>
<position>92,-23.5</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>GA_LED</type>
<position>75.5,-89</position>
<input>
<ID>N_in3</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_INVERTER</type>
<position>87.5,-84.5</position>
<input>
<ID>IN_0</ID>75 </input>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>121</ID>
<type>GA_LED</type>
<position>91.5,-84.5</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>DA_FROM</type>
<position>-10,-108</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>-8.5,-104</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_INVERTER</type>
<position>-2,-104</position>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_AND2</type>
<position>7,-106</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>GA_LED</type>
<position>13,-103</position>
<input>
<ID>N_in0</ID>86 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>DA_FROM</type>
<position>-8.5,-113.5</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>-10,-117.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_INVERTER</type>
<position>-1,-113.5</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_AND2</type>
<position>7,-115.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>13,-119</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>DA_FROM</type>
<position>-8.5,-100</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>133</ID>
<type>AI_XOR2</type>
<position>23,-105</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>86 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>GA_LED</type>
<position>27,-100.5</position>
<input>
<ID>N_in0</ID>87 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>DA_FROM</type>
<position>-8.5,-121.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>136</ID>
<type>AI_XOR2</type>
<position>22.5,-118.5</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>26.5,-121.5</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_AND2</type>
<position>36,-103.5</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>139</ID>
<type>GA_LED</type>
<position>41,-98</position>
<input>
<ID>N_in0</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_FULLADDER_1BIT</type>
<position>37,-115</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_B_0</ID>87 </input>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>141</ID>
<type>GA_LED</type>
<position>37,-122.5</position>
<input>
<ID>N_in3</ID>90 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>-10.5,-111</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_INVERTER</type>
<position>44,-108</position>
<input>
<ID>IN_0</ID>94 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND2</type>
<position>51.5,-100.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>51.5,-115.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AE_OR2</type>
<position>61,-107.5</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>91 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>55.5,-98.5</position>
<input>
<ID>N_in2</ID>96 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>55.5,-120.5</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>DA_FROM</type>
<position>-8.5,-96</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>150</ID>
<type>AI_XOR2</type>
<position>72,-107.5</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>65,-112</position>
<input>
<ID>N_in3</ID>92 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>78,-107.5</position>
<input>
<ID>N_in0</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>AE_OR2</type>
<position>78,-114</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>100 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>75.5,-118.5</position>
<input>
<ID>N_in3</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_INVERTER</type>
<position>87.5,-114</position>
<input>
<ID>IN_0</ID>98 </input>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>91.5,-114</position>
<input>
<ID>N_in0</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>-10,-138</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>158</ID>
<type>DA_FROM</type>
<position>-8.5,-134</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_INVERTER</type>
<position>-2,-134</position>
<input>
<ID>IN_0</ID>101 </input>
<output>
<ID>OUT_0</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_AND2</type>
<position>7,-136</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>GA_LED</type>
<position>13,-133</position>
<input>
<ID>N_in0</ID>109 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>DA_FROM</type>
<position>-8.5,-143.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>-10,-147.5</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_INVERTER</type>
<position>-1,-143.5</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_AND2</type>
<position>7,-145.5</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>GA_LED</type>
<position>13,-149</position>
<input>
<ID>N_in0</ID>107 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>-8.5,-130</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>168</ID>
<type>AI_XOR2</type>
<position>23,-135</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>27,-130.5</position>
<input>
<ID>N_in0</ID>110 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>DA_FROM</type>
<position>-8.5,-151.5</position>
<input>
<ID>IN_0</ID>111 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>171</ID>
<type>AI_XOR2</type>
<position>22.5,-148.5</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>111 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>GA_LED</type>
<position>26.5,-151.5</position>
<input>
<ID>N_in0</ID>112 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>36,-133.5</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>GA_LED</type>
<position>41,-128</position>
<input>
<ID>N_in0</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_FULLADDER_1BIT</type>
<position>37,-145</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_B_0</ID>110 </input>
<output>
<ID>OUT_0</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>176</ID>
<type>GA_LED</type>
<position>37,-152.5</position>
<input>
<ID>N_in3</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>DA_FROM</type>
<position>-10.5,-141</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_INVERTER</type>
<position>44,-138</position>
<input>
<ID>IN_0</ID>117 </input>
<output>
<ID>OUT_0</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND2</type>
<position>51.5,-130.5</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>118 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_AND2</type>
<position>51.5,-145.5</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>113 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>AE_OR2</type>
<position>61,-137.5</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>GA_LED</type>
<position>55.5,-128.5</position>
<input>
<ID>N_in2</ID>119 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>GA_LED</type>
<position>55.5,-150.5</position>
<input>
<ID>N_in0</ID>114 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>DA_FROM</type>
<position>-8.5,-126</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>185</ID>
<type>AI_XOR2</type>
<position>72,-137.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>GA_LED</type>
<position>65,-142</position>
<input>
<ID>N_in3</ID>115 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>GA_LED</type>
<position>78,-137.5</position>
<input>
<ID>N_in0</ID>123 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AE_OR2</type>
<position>78,-144</position>
<input>
<ID>IN_0</ID>123 </input>
<input>
<ID>IN_1</ID>123 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>GA_LED</type>
<position>75.5,-148.5</position>
<input>
<ID>N_in3</ID>123 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_INVERTER</type>
<position>87.5,-144</position>
<input>
<ID>IN_0</ID>121 </input>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>191</ID>
<type>GA_LED</type>
<position>91.5,-144</position>
<input>
<ID>N_in0</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>-10,-167.5</position>
<input>
<ID>IN_0</ID>126 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>193</ID>
<type>DA_FROM</type>
<position>-8.5,-163.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_INVERTER</type>
<position>-2,-163.5</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>195</ID>
<type>AA_AND2</type>
<position>7,-165.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>GA_LED</type>
<position>13,-162.5</position>
<input>
<ID>N_in0</ID>132 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>DA_FROM</type>
<position>-8.5,-173</position>
<input>
<ID>IN_0</ID>127 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>198</ID>
<type>DA_FROM</type>
<position>-10,-177</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_INVERTER</type>
<position>-1,-173</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND2</type>
<position>7,-175</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>GA_LED</type>
<position>13,-178.5</position>
<input>
<ID>N_in0</ID>130 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>-8.5,-159.5</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>203</ID>
<type>AI_XOR2</type>
<position>23,-164.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>132 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>GA_LED</type>
<position>27,-160</position>
<input>
<ID>N_in0</ID>133 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>DA_FROM</type>
<position>-8.5,-181</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>206</ID>
<type>AI_XOR2</type>
<position>22.5,-178</position>
<input>
<ID>IN_0</ID>130 </input>
<input>
<ID>IN_1</ID>134 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>GA_LED</type>
<position>26.5,-181</position>
<input>
<ID>N_in0</ID>135 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_AND2</type>
<position>36,-163</position>
<input>
<ID>IN_0</ID>133 </input>
<input>
<ID>IN_1</ID>135 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>209</ID>
<type>GA_LED</type>
<position>41,-157.5</position>
<input>
<ID>N_in0</ID>139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>210</ID>
<type>AA_FULLADDER_1BIT</type>
<position>37,-174.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_B_0</ID>133 </input>
<output>
<ID>OUT_0</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>211</ID>
<type>GA_LED</type>
<position>37,-182</position>
<input>
<ID>N_in3</ID>136 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>DA_FROM</type>
<position>-10.5,-170.5</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_INVERTER</type>
<position>44,-167.5</position>
<input>
<ID>IN_0</ID>140 </input>
<output>
<ID>OUT_0</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>51.5,-160</position>
<input>
<ID>IN_0</ID>139 </input>
<input>
<ID>IN_1</ID>141 </input>
<output>
<ID>OUT</ID>142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AA_AND2</type>
<position>51.5,-175</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>136 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AE_OR2</type>
<position>61,-167</position>
<input>
<ID>IN_0</ID>142 </input>
<input>
<ID>IN_1</ID>137 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>GA_LED</type>
<position>55.5,-158</position>
<input>
<ID>N_in2</ID>142 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>GA_LED</type>
<position>55.5,-180</position>
<input>
<ID>N_in0</ID>137 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>DA_FROM</type>
<position>-8.5,-155.5</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>220</ID>
<type>AI_XOR2</type>
<position>72,-167</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>138 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>GA_LED</type>
<position>65,-171.5</position>
<input>
<ID>N_in3</ID>138 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>GA_LED</type>
<position>78,-167</position>
<input>
<ID>N_in0</ID>146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AE_OR2</type>
<position>78,-173.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>146 </input>
<output>
<ID>OUT</ID>144 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>GA_LED</type>
<position>75.5,-178</position>
<input>
<ID>N_in3</ID>146 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>225</ID>
<type>AA_INVERTER</type>
<position>87.5,-173.5</position>
<input>
<ID>IN_0</ID>144 </input>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>226</ID>
<type>GA_LED</type>
<position>91.5,-173.5</position>
<input>
<ID>N_in0</ID>145 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>-12,-200.5</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>228</ID>
<type>DA_FROM</type>
<position>-10.5,-196.5</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_INVERTER</type>
<position>-4,-196.5</position>
<input>
<ID>IN_0</ID>147 </input>
<output>
<ID>OUT_0</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_AND2</type>
<position>5,-198.5</position>
<input>
<ID>IN_0</ID>148 </input>
<input>
<ID>IN_1</ID>149 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>231</ID>
<type>GA_LED</type>
<position>11,-195.5</position>
<input>
<ID>N_in0</ID>155 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>DA_FROM</type>
<position>-10.5,-206</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>233</ID>
<type>DA_FROM</type>
<position>-12,-210</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_INVERTER</type>
<position>-3,-206</position>
<input>
<ID>IN_0</ID>150 </input>
<output>
<ID>OUT_0</ID>151 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>235</ID>
<type>AA_AND2</type>
<position>5,-208</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>236</ID>
<type>GA_LED</type>
<position>11,-211.5</position>
<input>
<ID>N_in0</ID>153 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>237</ID>
<type>DA_FROM</type>
<position>-10.5,-192.5</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>238</ID>
<type>AI_XOR2</type>
<position>21,-197.5</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>155 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>GA_LED</type>
<position>25,-193</position>
<input>
<ID>N_in0</ID>156 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>240</ID>
<type>DA_FROM</type>
<position>-10.5,-214</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>241</ID>
<type>AI_XOR2</type>
<position>20.5,-211</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>242</ID>
<type>GA_LED</type>
<position>24.5,-214</position>
<input>
<ID>N_in0</ID>158 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>243</ID>
<type>AA_AND2</type>
<position>34,-196</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>158 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>GA_LED</type>
<position>39,-190.5</position>
<input>
<ID>N_in0</ID>162 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>245</ID>
<type>AA_FULLADDER_1BIT</type>
<position>35,-207.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_B_0</ID>156 </input>
<output>
<ID>OUT_0</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>246</ID>
<type>GA_LED</type>
<position>35,-215</position>
<input>
<ID>N_in3</ID>159 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>DA_FROM</type>
<position>-12.5,-203.5</position>
<input>
<ID>IN_0</ID>163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>248</ID>
<type>AA_INVERTER</type>
<position>42,-200.5</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>249</ID>
<type>AA_AND2</type>
<position>49.5,-193</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>164 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_AND2</type>
<position>49.5,-208</position>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>AE_OR2</type>
<position>59,-200</position>
<input>
<ID>IN_0</ID>165 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>252</ID>
<type>GA_LED</type>
<position>53.5,-191</position>
<input>
<ID>N_in2</ID>165 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>GA_LED</type>
<position>53.5,-213</position>
<input>
<ID>N_in0</ID>160 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>254</ID>
<type>DA_FROM</type>
<position>-10.5,-188.5</position>
<input>
<ID>IN_0</ID>166 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>255</ID>
<type>AI_XOR2</type>
<position>70,-200</position>
<input>
<ID>IN_0</ID>166 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>GA_LED</type>
<position>63,-204.5</position>
<input>
<ID>N_in3</ID>161 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>257</ID>
<type>GA_LED</type>
<position>76,-200</position>
<input>
<ID>N_in0</ID>169 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>AE_OR2</type>
<position>76,-206.5</position>
<input>
<ID>IN_0</ID>169 </input>
<input>
<ID>IN_1</ID>169 </input>
<output>
<ID>OUT</ID>167 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>259</ID>
<type>GA_LED</type>
<position>73.5,-211</position>
<input>
<ID>N_in3</ID>169 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>260</ID>
<type>AA_INVERTER</type>
<position>85.5,-206.5</position>
<input>
<ID>IN_0</ID>167 </input>
<output>
<ID>OUT_0</ID>168 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>261</ID>
<type>GA_LED</type>
<position>89.5,-206.5</position>
<input>
<ID>N_in0</ID>168 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>DA_FROM</type>
<position>130,-19.5</position>
<input>
<ID>IN_0</ID>172 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>263</ID>
<type>DA_FROM</type>
<position>131.5,-15.5</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_INVERTER</type>
<position>138,-15.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>171 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>265</ID>
<type>AA_AND2</type>
<position>147,-17.5</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>266</ID>
<type>GA_LED</type>
<position>153,-14.5</position>
<input>
<ID>N_in0</ID>178 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>DA_FROM</type>
<position>131.5,-25</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>268</ID>
<type>DA_FROM</type>
<position>130,-29</position>
<input>
<ID>IN_0</ID>175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>269</ID>
<type>AA_INVERTER</type>
<position>139,-25</position>
<input>
<ID>IN_0</ID>173 </input>
<output>
<ID>OUT_0</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>270</ID>
<type>AA_AND2</type>
<position>147,-27</position>
<input>
<ID>IN_0</ID>174 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>271</ID>
<type>GA_LED</type>
<position>153,-30.5</position>
<input>
<ID>N_in0</ID>176 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>272</ID>
<type>DA_FROM</type>
<position>131.5,-11.5</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>273</ID>
<type>AI_XOR2</type>
<position>163,-16.5</position>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>274</ID>
<type>GA_LED</type>
<position>167,-12</position>
<input>
<ID>N_in0</ID>179 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>275</ID>
<type>DA_FROM</type>
<position>131.5,-33</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>276</ID>
<type>AI_XOR2</type>
<position>162.5,-30</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>180 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>GA_LED</type>
<position>166.5,-33</position>
<input>
<ID>N_in0</ID>181 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>176,-15</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>GA_LED</type>
<position>181,-9.5</position>
<input>
<ID>N_in0</ID>185 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>280</ID>
<type>AA_FULLADDER_1BIT</type>
<position>177,-26.5</position>
<input>
<ID>IN_0</ID>181 </input>
<input>
<ID>IN_B_0</ID>179 </input>
<output>
<ID>OUT_0</ID>182 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>281</ID>
<type>GA_LED</type>
<position>177,-34</position>
<input>
<ID>N_in3</ID>182 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>282</ID>
<type>DA_FROM</type>
<position>129.5,-22.5</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>283</ID>
<type>AA_INVERTER</type>
<position>184,-19.5</position>
<input>
<ID>IN_0</ID>186 </input>
<output>
<ID>OUT_0</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>284</ID>
<type>AA_AND2</type>
<position>191.5,-12</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>285</ID>
<type>AA_AND2</type>
<position>191.5,-27</position>
<input>
<ID>IN_0</ID>186 </input>
<input>
<ID>IN_1</ID>182 </input>
<output>
<ID>OUT</ID>183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>AE_OR2</type>
<position>201,-19</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>183 </input>
<output>
<ID>OUT</ID>184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>287</ID>
<type>GA_LED</type>
<position>195.5,-10</position>
<input>
<ID>N_in2</ID>188 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>288</ID>
<type>GA_LED</type>
<position>195.5,-32</position>
<input>
<ID>N_in0</ID>183 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>DA_FROM</type>
<position>131.5,-7.5</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>290</ID>
<type>AI_XOR2</type>
<position>212,-19</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>291</ID>
<type>GA_LED</type>
<position>205,-23.5</position>
<input>
<ID>N_in3</ID>184 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>292</ID>
<type>GA_LED</type>
<position>218,-19</position>
<input>
<ID>N_in0</ID>192 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AE_OR2</type>
<position>218,-25.5</position>
<input>
<ID>IN_0</ID>192 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>190 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>294</ID>
<type>GA_LED</type>
<position>215.5,-30</position>
<input>
<ID>N_in3</ID>192 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>295</ID>
<type>AA_INVERTER</type>
<position>227.5,-25.5</position>
<input>
<ID>IN_0</ID>190 </input>
<output>
<ID>OUT_0</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>296</ID>
<type>GA_LED</type>
<position>231.5,-25.5</position>
<input>
<ID>N_in0</ID>191 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>297</ID>
<type>DA_FROM</type>
<position>130,-50.5</position>
<input>
<ID>IN_0</ID>195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>298</ID>
<type>DA_FROM</type>
<position>131.5,-46.5</position>
<input>
<ID>IN_0</ID>193 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_INVERTER</type>
<position>138,-46.5</position>
<input>
<ID>IN_0</ID>193 </input>
<output>
<ID>OUT_0</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_AND2</type>
<position>147,-48.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>195 </input>
<output>
<ID>OUT</ID>201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>GA_LED</type>
<position>153,-45.5</position>
<input>
<ID>N_in0</ID>201 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>302</ID>
<type>DA_FROM</type>
<position>131.5,-56</position>
<input>
<ID>IN_0</ID>196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>303</ID>
<type>DA_FROM</type>
<position>130,-60</position>
<input>
<ID>IN_0</ID>198 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_INVERTER</type>
<position>139,-56</position>
<input>
<ID>IN_0</ID>196 </input>
<output>
<ID>OUT_0</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>305</ID>
<type>AA_AND2</type>
<position>147,-58</position>
<input>
<ID>IN_0</ID>197 </input>
<input>
<ID>IN_1</ID>198 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>306</ID>
<type>GA_LED</type>
<position>153,-61.5</position>
<input>
<ID>N_in0</ID>199 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>131.5,-42.5</position>
<input>
<ID>IN_0</ID>200 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>308</ID>
<type>AI_XOR2</type>
<position>163,-47.5</position>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>201 </input>
<output>
<ID>OUT</ID>202 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>GA_LED</type>
<position>167,-43</position>
<input>
<ID>N_in0</ID>202 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>DA_FROM</type>
<position>131.5,-64</position>
<input>
<ID>IN_0</ID>203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>311</ID>
<type>AI_XOR2</type>
<position>162.5,-61</position>
<input>
<ID>IN_0</ID>199 </input>
<input>
<ID>IN_1</ID>203 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>312</ID>
<type>GA_LED</type>
<position>166.5,-64</position>
<input>
<ID>N_in0</ID>204 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>313</ID>
<type>AA_AND2</type>
<position>176,-46</position>
<input>
<ID>IN_0</ID>202 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>208 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>314</ID>
<type>GA_LED</type>
<position>181,-40.5</position>
<input>
<ID>N_in0</ID>208 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>315</ID>
<type>AA_FULLADDER_1BIT</type>
<position>177,-57.5</position>
<input>
<ID>IN_0</ID>204 </input>
<input>
<ID>IN_B_0</ID>202 </input>
<output>
<ID>OUT_0</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>316</ID>
<type>GA_LED</type>
<position>177,-65</position>
<input>
<ID>N_in3</ID>205 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>129.5,-53.5</position>
<input>
<ID>IN_0</ID>209 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_INVERTER</type>
<position>184,-50.5</position>
<input>
<ID>IN_0</ID>209 </input>
<output>
<ID>OUT_0</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_AND2</type>
<position>191.5,-43</position>
<input>
<ID>IN_0</ID>208 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>320</ID>
<type>AA_AND2</type>
<position>191.5,-58</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>AE_OR2</type>
<position>201,-50</position>
<input>
<ID>IN_0</ID>211 </input>
<input>
<ID>IN_1</ID>206 </input>
<output>
<ID>OUT</ID>207 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>322</ID>
<type>GA_LED</type>
<position>195.5,-41</position>
<input>
<ID>N_in2</ID>211 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>323</ID>
<type>GA_LED</type>
<position>195.5,-63</position>
<input>
<ID>N_in0</ID>206 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>324</ID>
<type>DA_FROM</type>
<position>131.5,-38.5</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>325</ID>
<type>AI_XOR2</type>
<position>212,-50</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>207 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>326</ID>
<type>GA_LED</type>
<position>205,-54.5</position>
<input>
<ID>N_in3</ID>207 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>327</ID>
<type>GA_LED</type>
<position>218,-50</position>
<input>
<ID>N_in0</ID>215 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>328</ID>
<type>AE_OR2</type>
<position>218,-56.5</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>215 </input>
<output>
<ID>OUT</ID>213 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>GA_LED</type>
<position>215.5,-61</position>
<input>
<ID>N_in3</ID>215 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>330</ID>
<type>AA_INVERTER</type>
<position>227.5,-56.5</position>
<input>
<ID>IN_0</ID>213 </input>
<output>
<ID>OUT_0</ID>214 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>331</ID>
<type>GA_LED</type>
<position>231.5,-56.5</position>
<input>
<ID>N_in0</ID>214 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>332</ID>
<type>DA_FROM</type>
<position>131,-82.5</position>
<input>
<ID>IN_0</ID>218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>132.5,-78.5</position>
<input>
<ID>IN_0</ID>216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>334</ID>
<type>AA_INVERTER</type>
<position>139,-78.5</position>
<input>
<ID>IN_0</ID>216 </input>
<output>
<ID>OUT_0</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>335</ID>
<type>AA_AND2</type>
<position>148,-80.5</position>
<input>
<ID>IN_0</ID>217 </input>
<input>
<ID>IN_1</ID>218 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>336</ID>
<type>GA_LED</type>
<position>154,-77.5</position>
<input>
<ID>N_in0</ID>224 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>337</ID>
<type>DA_FROM</type>
<position>132.5,-88</position>
<input>
<ID>IN_0</ID>219 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>338</ID>
<type>DA_FROM</type>
<position>131,-92</position>
<input>
<ID>IN_0</ID>221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>339</ID>
<type>AA_INVERTER</type>
<position>140,-88</position>
<input>
<ID>IN_0</ID>219 </input>
<output>
<ID>OUT_0</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_AND2</type>
<position>148,-90</position>
<input>
<ID>IN_0</ID>220 </input>
<input>
<ID>IN_1</ID>221 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>GA_LED</type>
<position>154,-93.5</position>
<input>
<ID>N_in0</ID>222 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>342</ID>
<type>DA_FROM</type>
<position>132.5,-74.5</position>
<input>
<ID>IN_0</ID>223 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>343</ID>
<type>AI_XOR2</type>
<position>164,-79.5</position>
<input>
<ID>IN_0</ID>223 </input>
<input>
<ID>IN_1</ID>224 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>344</ID>
<type>GA_LED</type>
<position>168,-75</position>
<input>
<ID>N_in0</ID>225 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>345</ID>
<type>DA_FROM</type>
<position>132.5,-96</position>
<input>
<ID>IN_0</ID>226 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>346</ID>
<type>AI_XOR2</type>
<position>163.5,-93</position>
<input>
<ID>IN_0</ID>222 </input>
<input>
<ID>IN_1</ID>226 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>347</ID>
<type>GA_LED</type>
<position>167.5,-96</position>
<input>
<ID>N_in0</ID>227 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>348</ID>
<type>AA_AND2</type>
<position>177,-78</position>
<input>
<ID>IN_0</ID>225 </input>
<input>
<ID>IN_1</ID>227 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>GA_LED</type>
<position>182,-72.5</position>
<input>
<ID>N_in0</ID>231 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>AA_FULLADDER_1BIT</type>
<position>178,-89.5</position>
<input>
<ID>IN_0</ID>227 </input>
<input>
<ID>IN_B_0</ID>225 </input>
<output>
<ID>OUT_0</ID>228 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>351</ID>
<type>GA_LED</type>
<position>178,-97</position>
<input>
<ID>N_in3</ID>228 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>352</ID>
<type>DA_FROM</type>
<position>130.5,-85.5</position>
<input>
<ID>IN_0</ID>232 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>353</ID>
<type>AA_INVERTER</type>
<position>185,-82.5</position>
<input>
<ID>IN_0</ID>232 </input>
<output>
<ID>OUT_0</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_AND2</type>
<position>192.5,-75</position>
<input>
<ID>IN_0</ID>231 </input>
<input>
<ID>IN_1</ID>233 </input>
<output>
<ID>OUT</ID>234 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_AND2</type>
<position>192.5,-90</position>
<input>
<ID>IN_0</ID>232 </input>
<input>
<ID>IN_1</ID>228 </input>
<output>
<ID>OUT</ID>229 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>356</ID>
<type>AE_OR2</type>
<position>202,-82</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>229 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>GA_LED</type>
<position>196.5,-73</position>
<input>
<ID>N_in2</ID>234 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>358</ID>
<type>GA_LED</type>
<position>196.5,-95</position>
<input>
<ID>N_in0</ID>229 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>359</ID>
<type>DA_FROM</type>
<position>132.5,-70.5</position>
<input>
<ID>IN_0</ID>235 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>360</ID>
<type>AI_XOR2</type>
<position>213,-82</position>
<input>
<ID>IN_0</ID>235 </input>
<input>
<ID>IN_1</ID>230 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>GA_LED</type>
<position>206,-86.5</position>
<input>
<ID>N_in3</ID>230 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>362</ID>
<type>GA_LED</type>
<position>219,-82</position>
<input>
<ID>N_in0</ID>238 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>363</ID>
<type>AE_OR2</type>
<position>219,-88.5</position>
<input>
<ID>IN_0</ID>238 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>364</ID>
<type>GA_LED</type>
<position>216.5,-93</position>
<input>
<ID>N_in3</ID>238 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>365</ID>
<type>AA_INVERTER</type>
<position>228.5,-88.5</position>
<input>
<ID>IN_0</ID>236 </input>
<output>
<ID>OUT_0</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>366</ID>
<type>GA_LED</type>
<position>232.5,-88.5</position>
<input>
<ID>N_in0</ID>237 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>367</ID>
<type>DA_FROM</type>
<position>132,-113.5</position>
<input>
<ID>IN_0</ID>241 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>368</ID>
<type>DA_FROM</type>
<position>133.5,-109.5</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_INVERTER</type>
<position>140,-109.5</position>
<input>
<ID>IN_0</ID>239 </input>
<output>
<ID>OUT_0</ID>240 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>370</ID>
<type>AA_AND2</type>
<position>149,-111.5</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>371</ID>
<type>GA_LED</type>
<position>155,-108.5</position>
<input>
<ID>N_in0</ID>247 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>372</ID>
<type>DA_FROM</type>
<position>133.5,-119</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>373</ID>
<type>DA_FROM</type>
<position>132,-123</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>374</ID>
<type>AA_INVERTER</type>
<position>141,-119</position>
<input>
<ID>IN_0</ID>242 </input>
<output>
<ID>OUT_0</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>375</ID>
<type>AA_AND2</type>
<position>149,-121</position>
<input>
<ID>IN_0</ID>243 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>376</ID>
<type>GA_LED</type>
<position>155,-124.5</position>
<input>
<ID>N_in0</ID>245 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>377</ID>
<type>DA_FROM</type>
<position>133.5,-105.5</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>378</ID>
<type>AI_XOR2</type>
<position>165,-110.5</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>247 </input>
<output>
<ID>OUT</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>379</ID>
<type>GA_LED</type>
<position>169,-106</position>
<input>
<ID>N_in0</ID>248 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>380</ID>
<type>DA_FROM</type>
<position>133.5,-127</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>381</ID>
<type>AI_XOR2</type>
<position>164.5,-124</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>249 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>382</ID>
<type>GA_LED</type>
<position>168.5,-127</position>
<input>
<ID>N_in0</ID>250 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>383</ID>
<type>AA_AND2</type>
<position>178,-109</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>GA_LED</type>
<position>183,-103.5</position>
<input>
<ID>N_in0</ID>254 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>385</ID>
<type>AA_FULLADDER_1BIT</type>
<position>179,-120.5</position>
<input>
<ID>IN_0</ID>250 </input>
<input>
<ID>IN_B_0</ID>248 </input>
<output>
<ID>OUT_0</ID>251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>386</ID>
<type>GA_LED</type>
<position>179,-128</position>
<input>
<ID>N_in3</ID>251 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>387</ID>
<type>DA_FROM</type>
<position>131.5,-116.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>388</ID>
<type>AA_INVERTER</type>
<position>186,-113.5</position>
<input>
<ID>IN_0</ID>255 </input>
<output>
<ID>OUT_0</ID>256 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>389</ID>
<type>AA_AND2</type>
<position>193.5,-106</position>
<input>
<ID>IN_0</ID>254 </input>
<input>
<ID>IN_1</ID>256 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>390</ID>
<type>AA_AND2</type>
<position>193.5,-121</position>
<input>
<ID>IN_0</ID>255 </input>
<input>
<ID>IN_1</ID>251 </input>
<output>
<ID>OUT</ID>252 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>391</ID>
<type>AE_OR2</type>
<position>203,-113</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>252 </input>
<output>
<ID>OUT</ID>253 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>392</ID>
<type>GA_LED</type>
<position>197.5,-104</position>
<input>
<ID>N_in2</ID>257 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>393</ID>
<type>GA_LED</type>
<position>197.5,-126</position>
<input>
<ID>N_in0</ID>252 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>394</ID>
<type>DA_FROM</type>
<position>133.5,-101.5</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>395</ID>
<type>AI_XOR2</type>
<position>214,-113</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>396</ID>
<type>GA_LED</type>
<position>207,-117.5</position>
<input>
<ID>N_in3</ID>253 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>397</ID>
<type>GA_LED</type>
<position>220,-113</position>
<input>
<ID>N_in0</ID>261 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>398</ID>
<type>AE_OR2</type>
<position>220,-119.5</position>
<input>
<ID>IN_0</ID>261 </input>
<input>
<ID>IN_1</ID>261 </input>
<output>
<ID>OUT</ID>259 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>399</ID>
<type>GA_LED</type>
<position>217.5,-124</position>
<input>
<ID>N_in3</ID>261 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>400</ID>
<type>AA_INVERTER</type>
<position>229.5,-119.5</position>
<input>
<ID>IN_0</ID>259 </input>
<output>
<ID>OUT_0</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>401</ID>
<type>GA_LED</type>
<position>233.5,-119.5</position>
<input>
<ID>N_in0</ID>260 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>402</ID>
<type>DA_FROM</type>
<position>132,-144.5</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>403</ID>
<type>DA_FROM</type>
<position>133.5,-140.5</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_INVERTER</type>
<position>140,-140.5</position>
<input>
<ID>IN_0</ID>262 </input>
<output>
<ID>OUT_0</ID>263 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>405</ID>
<type>AA_AND2</type>
<position>149,-142.5</position>
<input>
<ID>IN_0</ID>263 </input>
<input>
<ID>IN_1</ID>264 </input>
<output>
<ID>OUT</ID>270 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>406</ID>
<type>GA_LED</type>
<position>155,-139.5</position>
<input>
<ID>N_in0</ID>270 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>407</ID>
<type>DA_FROM</type>
<position>133.5,-150</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>408</ID>
<type>DA_FROM</type>
<position>132,-154</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_INVERTER</type>
<position>141,-150</position>
<input>
<ID>IN_0</ID>265 </input>
<output>
<ID>OUT_0</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>410</ID>
<type>AA_AND2</type>
<position>149,-152</position>
<input>
<ID>IN_0</ID>266 </input>
<input>
<ID>IN_1</ID>267 </input>
<output>
<ID>OUT</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>411</ID>
<type>GA_LED</type>
<position>155,-155.5</position>
<input>
<ID>N_in0</ID>268 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>133.5,-136.5</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>413</ID>
<type>AI_XOR2</type>
<position>165,-141.5</position>
<input>
<ID>IN_0</ID>269 </input>
<input>
<ID>IN_1</ID>270 </input>
<output>
<ID>OUT</ID>271 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>414</ID>
<type>GA_LED</type>
<position>169,-137</position>
<input>
<ID>N_in0</ID>271 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>415</ID>
<type>DA_FROM</type>
<position>133.5,-158</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>416</ID>
<type>AI_XOR2</type>
<position>164.5,-155</position>
<input>
<ID>IN_0</ID>268 </input>
<input>
<ID>IN_1</ID>272 </input>
<output>
<ID>OUT</ID>273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>GA_LED</type>
<position>168.5,-158</position>
<input>
<ID>N_in0</ID>273 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>418</ID>
<type>AA_AND2</type>
<position>178,-140</position>
<input>
<ID>IN_0</ID>271 </input>
<input>
<ID>IN_1</ID>273 </input>
<output>
<ID>OUT</ID>277 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>419</ID>
<type>GA_LED</type>
<position>183,-134.5</position>
<input>
<ID>N_in0</ID>277 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>420</ID>
<type>AA_FULLADDER_1BIT</type>
<position>179,-151.5</position>
<input>
<ID>IN_0</ID>273 </input>
<input>
<ID>IN_B_0</ID>271 </input>
<output>
<ID>OUT_0</ID>274 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>421</ID>
<type>GA_LED</type>
<position>179,-159</position>
<input>
<ID>N_in3</ID>274 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>422</ID>
<type>DA_FROM</type>
<position>131.5,-147.5</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>423</ID>
<type>AA_INVERTER</type>
<position>186,-144.5</position>
<input>
<ID>IN_0</ID>278 </input>
<output>
<ID>OUT_0</ID>279 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>424</ID>
<type>AA_AND2</type>
<position>193.5,-137</position>
<input>
<ID>IN_0</ID>277 </input>
<input>
<ID>IN_1</ID>279 </input>
<output>
<ID>OUT</ID>280 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>425</ID>
<type>AA_AND2</type>
<position>193.5,-152</position>
<input>
<ID>IN_0</ID>278 </input>
<input>
<ID>IN_1</ID>274 </input>
<output>
<ID>OUT</ID>275 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>426</ID>
<type>AE_OR2</type>
<position>203,-144</position>
<input>
<ID>IN_0</ID>280 </input>
<input>
<ID>IN_1</ID>275 </input>
<output>
<ID>OUT</ID>276 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>427</ID>
<type>GA_LED</type>
<position>197.5,-135</position>
<input>
<ID>N_in2</ID>280 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>428</ID>
<type>GA_LED</type>
<position>197.5,-157</position>
<input>
<ID>N_in0</ID>275 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>429</ID>
<type>DA_FROM</type>
<position>133.5,-132.5</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>430</ID>
<type>AI_XOR2</type>
<position>214,-144</position>
<input>
<ID>IN_0</ID>281 </input>
<input>
<ID>IN_1</ID>276 </input>
<output>
<ID>OUT</ID>284 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>431</ID>
<type>GA_LED</type>
<position>207,-148.5</position>
<input>
<ID>N_in3</ID>276 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>432</ID>
<type>GA_LED</type>
<position>220,-144</position>
<input>
<ID>N_in0</ID>284 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>433</ID>
<type>AE_OR2</type>
<position>220,-150.5</position>
<input>
<ID>IN_0</ID>284 </input>
<input>
<ID>IN_1</ID>284 </input>
<output>
<ID>OUT</ID>282 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>434</ID>
<type>GA_LED</type>
<position>217.5,-155</position>
<input>
<ID>N_in3</ID>284 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>435</ID>
<type>AA_INVERTER</type>
<position>229.5,-150.5</position>
<input>
<ID>IN_0</ID>282 </input>
<output>
<ID>OUT_0</ID>283 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>436</ID>
<type>GA_LED</type>
<position>233.5,-150.5</position>
<input>
<ID>N_in0</ID>283 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>437</ID>
<type>DA_FROM</type>
<position>130,-174.5</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>438</ID>
<type>DA_FROM</type>
<position>131.5,-170.5</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>439</ID>
<type>AA_INVERTER</type>
<position>138,-170.5</position>
<input>
<ID>IN_0</ID>285 </input>
<output>
<ID>OUT_0</ID>286 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>440</ID>
<type>AA_AND2</type>
<position>147,-172.5</position>
<input>
<ID>IN_0</ID>286 </input>
<input>
<ID>IN_1</ID>287 </input>
<output>
<ID>OUT</ID>293 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>441</ID>
<type>GA_LED</type>
<position>153,-169.5</position>
<input>
<ID>N_in0</ID>293 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>442</ID>
<type>DA_FROM</type>
<position>131.5,-180</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>443</ID>
<type>DA_FROM</type>
<position>130,-184</position>
<input>
<ID>IN_0</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>444</ID>
<type>AA_INVERTER</type>
<position>139,-180</position>
<input>
<ID>IN_0</ID>288 </input>
<output>
<ID>OUT_0</ID>289 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>445</ID>
<type>AA_AND2</type>
<position>147,-182</position>
<input>
<ID>IN_0</ID>289 </input>
<input>
<ID>IN_1</ID>290 </input>
<output>
<ID>OUT</ID>291 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>446</ID>
<type>GA_LED</type>
<position>153,-185.5</position>
<input>
<ID>N_in0</ID>291 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>131.5,-166.5</position>
<input>
<ID>IN_0</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>448</ID>
<type>AI_XOR2</type>
<position>163,-171.5</position>
<input>
<ID>IN_0</ID>292 </input>
<input>
<ID>IN_1</ID>293 </input>
<output>
<ID>OUT</ID>294 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>449</ID>
<type>GA_LED</type>
<position>167,-167</position>
<input>
<ID>N_in0</ID>294 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>450</ID>
<type>DA_FROM</type>
<position>131.5,-188</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>451</ID>
<type>AI_XOR2</type>
<position>162.5,-185</position>
<input>
<ID>IN_0</ID>291 </input>
<input>
<ID>IN_1</ID>295 </input>
<output>
<ID>OUT</ID>296 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>452</ID>
<type>GA_LED</type>
<position>166.5,-188</position>
<input>
<ID>N_in0</ID>296 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>453</ID>
<type>AA_AND2</type>
<position>176,-170</position>
<input>
<ID>IN_0</ID>294 </input>
<input>
<ID>IN_1</ID>296 </input>
<output>
<ID>OUT</ID>300 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>454</ID>
<type>GA_LED</type>
<position>181,-164.5</position>
<input>
<ID>N_in0</ID>300 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>455</ID>
<type>AA_FULLADDER_1BIT</type>
<position>177,-181.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_B_0</ID>294 </input>
<output>
<ID>OUT_0</ID>297 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>456</ID>
<type>GA_LED</type>
<position>177,-189</position>
<input>
<ID>N_in3</ID>297 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>457</ID>
<type>DA_FROM</type>
<position>129.5,-177.5</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>458</ID>
<type>AA_INVERTER</type>
<position>184,-174.5</position>
<input>
<ID>IN_0</ID>301 </input>
<output>
<ID>OUT_0</ID>302 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>459</ID>
<type>AA_AND2</type>
<position>191.5,-167</position>
<input>
<ID>IN_0</ID>300 </input>
<input>
<ID>IN_1</ID>302 </input>
<output>
<ID>OUT</ID>303 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>460</ID>
<type>AA_AND2</type>
<position>191.5,-182</position>
<input>
<ID>IN_0</ID>301 </input>
<input>
<ID>IN_1</ID>297 </input>
<output>
<ID>OUT</ID>298 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>461</ID>
<type>AE_OR2</type>
<position>201,-174</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>298 </input>
<output>
<ID>OUT</ID>299 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>462</ID>
<type>GA_LED</type>
<position>195.5,-165</position>
<input>
<ID>N_in2</ID>303 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>463</ID>
<type>GA_LED</type>
<position>195.5,-187</position>
<input>
<ID>N_in0</ID>298 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>464</ID>
<type>DA_FROM</type>
<position>131.5,-162.5</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>465</ID>
<type>AI_XOR2</type>
<position>212,-174</position>
<input>
<ID>IN_0</ID>304 </input>
<input>
<ID>IN_1</ID>299 </input>
<output>
<ID>OUT</ID>307 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>466</ID>
<type>GA_LED</type>
<position>205,-178.5</position>
<input>
<ID>N_in3</ID>299 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>467</ID>
<type>GA_LED</type>
<position>218,-174</position>
<input>
<ID>N_in0</ID>307 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>468</ID>
<type>AE_OR2</type>
<position>218,-180.5</position>
<input>
<ID>IN_0</ID>307 </input>
<input>
<ID>IN_1</ID>307 </input>
<output>
<ID>OUT</ID>305 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>469</ID>
<type>GA_LED</type>
<position>215.5,-185</position>
<input>
<ID>N_in3</ID>307 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>470</ID>
<type>AA_INVERTER</type>
<position>227.5,-180.5</position>
<input>
<ID>IN_0</ID>305 </input>
<output>
<ID>OUT_0</ID>306 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>471</ID>
<type>GA_LED</type>
<position>231.5,-180.5</position>
<input>
<ID>N_in0</ID>306 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>472</ID>
<type>DA_FROM</type>
<position>129,-206.5</position>
<input>
<ID>IN_0</ID>310 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID X</lparam></gate>
<gate>
<ID>473</ID>
<type>DA_FROM</type>
<position>130.5,-202.5</position>
<input>
<ID>IN_0</ID>308 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZX</lparam></gate>
<gate>
<ID>474</ID>
<type>AA_INVERTER</type>
<position>137,-202.5</position>
<input>
<ID>IN_0</ID>308 </input>
<output>
<ID>OUT_0</ID>309 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>475</ID>
<type>AA_AND2</type>
<position>146,-204.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>310 </input>
<output>
<ID>OUT</ID>316 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>476</ID>
<type>GA_LED</type>
<position>152,-201.5</position>
<input>
<ID>N_in0</ID>316 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>477</ID>
<type>DA_FROM</type>
<position>130.5,-212</position>
<input>
<ID>IN_0</ID>311 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ZY</lparam></gate>
<gate>
<ID>478</ID>
<type>DA_FROM</type>
<position>129,-216</position>
<input>
<ID>IN_0</ID>313 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Y</lparam></gate>
<gate>
<ID>479</ID>
<type>AA_INVERTER</type>
<position>138,-212</position>
<input>
<ID>IN_0</ID>311 </input>
<output>
<ID>OUT_0</ID>312 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>480</ID>
<type>AA_AND2</type>
<position>146,-214</position>
<input>
<ID>IN_0</ID>312 </input>
<input>
<ID>IN_1</ID>313 </input>
<output>
<ID>OUT</ID>314 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>481</ID>
<type>GA_LED</type>
<position>152,-217.5</position>
<input>
<ID>N_in0</ID>314 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>482</ID>
<type>DA_FROM</type>
<position>130.5,-198.5</position>
<input>
<ID>IN_0</ID>315 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NX</lparam></gate>
<gate>
<ID>483</ID>
<type>AI_XOR2</type>
<position>162,-203.5</position>
<input>
<ID>IN_0</ID>315 </input>
<input>
<ID>IN_1</ID>316 </input>
<output>
<ID>OUT</ID>317 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>484</ID>
<type>GA_LED</type>
<position>166,-199</position>
<input>
<ID>N_in0</ID>317 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>485</ID>
<type>DA_FROM</type>
<position>130.5,-220</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NY</lparam></gate>
<gate>
<ID>486</ID>
<type>AI_XOR2</type>
<position>161.5,-217</position>
<input>
<ID>IN_0</ID>314 </input>
<input>
<ID>IN_1</ID>318 </input>
<output>
<ID>OUT</ID>319 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>487</ID>
<type>GA_LED</type>
<position>165.5,-220</position>
<input>
<ID>N_in0</ID>319 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>488</ID>
<type>AA_AND2</type>
<position>175,-202</position>
<input>
<ID>IN_0</ID>317 </input>
<input>
<ID>IN_1</ID>319 </input>
<output>
<ID>OUT</ID>323 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>489</ID>
<type>GA_LED</type>
<position>180,-196.5</position>
<input>
<ID>N_in0</ID>323 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>490</ID>
<type>AA_FULLADDER_1BIT</type>
<position>176,-213.5</position>
<input>
<ID>IN_0</ID>319 </input>
<input>
<ID>IN_B_0</ID>317 </input>
<output>
<ID>OUT_0</ID>320 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>491</ID>
<type>GA_LED</type>
<position>176,-221</position>
<input>
<ID>N_in3</ID>320 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>492</ID>
<type>DA_FROM</type>
<position>128.5,-209.5</position>
<input>
<ID>IN_0</ID>324 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>493</ID>
<type>AA_INVERTER</type>
<position>183,-206.5</position>
<input>
<ID>IN_0</ID>324 </input>
<output>
<ID>OUT_0</ID>325 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_AND2</type>
<position>190.5,-199</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>325 </input>
<output>
<ID>OUT</ID>326 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>495</ID>
<type>AA_AND2</type>
<position>190.5,-214</position>
<input>
<ID>IN_0</ID>324 </input>
<input>
<ID>IN_1</ID>320 </input>
<output>
<ID>OUT</ID>321 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>496</ID>
<type>AE_OR2</type>
<position>200,-206</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>321 </input>
<output>
<ID>OUT</ID>322 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>497</ID>
<type>GA_LED</type>
<position>194.5,-197</position>
<input>
<ID>N_in2</ID>326 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>498</ID>
<type>GA_LED</type>
<position>194.5,-219</position>
<input>
<ID>N_in0</ID>321 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>499</ID>
<type>DA_FROM</type>
<position>130.5,-194.5</position>
<input>
<ID>IN_0</ID>327 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID NO</lparam></gate>
<gate>
<ID>500</ID>
<type>AI_XOR2</type>
<position>211,-206</position>
<input>
<ID>IN_0</ID>327 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>330 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>501</ID>
<type>GA_LED</type>
<position>204,-210.5</position>
<input>
<ID>N_in3</ID>322 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>502</ID>
<type>GA_LED</type>
<position>217,-206</position>
<input>
<ID>N_in0</ID>330 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>503</ID>
<type>AE_OR2</type>
<position>217,-212.5</position>
<input>
<ID>IN_0</ID>330 </input>
<input>
<ID>IN_1</ID>330 </input>
<output>
<ID>OUT</ID>328 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>504</ID>
<type>GA_LED</type>
<position>214.5,-217</position>
<input>
<ID>N_in3</ID>330 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>505</ID>
<type>AA_INVERTER</type>
<position>226.5,-212.5</position>
<input>
<ID>IN_0</ID>328 </input>
<output>
<ID>OUT_0</ID>329 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>506</ID>
<type>GA_LED</type>
<position>230.5,-212.5</position>
<input>
<ID>N_in0</ID>329 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-7,19,-6,19</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-7,15.5,-6,15.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<connection>
<GID>8</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-44.5,-4.5,-44.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-45.5,2.5,-44.5</points>
<intersection>-45.5 1</intersection>
<intersection>-44.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-45.5,4.5,-45.5</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-44.5,2.5,-44.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-48.5,-3,-47.5</points>
<intersection>-48.5 2</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3,-47.5,4.5,-47.5</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>-3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-48.5,-3,-48.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>-3 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-13.5,-4.5,-13.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-14.5,2.5,-13.5</points>
<intersection>-14.5 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-14.5,4.5,-14.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-13.5,2.5,-13.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-17.5,-3,-16.5</points>
<intersection>-17.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3,-16.5,4.5,-16.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-17.5,-3,-17.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-3 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-54,-3.5,-54</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,19,7,19</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7,12,-6,12</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6,-23,-3.5,-23</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-24,3.5,-23</points>
<intersection>-24 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-24,4.5,-24</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-23,3.5,-23</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-27,-0.5,-26</points>
<intersection>-27 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-26,4.5,-26</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-27,-0.5,-27</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-28.5,15,-25</points>
<intersection>-28.5 9</intersection>
<intersection>-27 10</intersection>
<intersection>-25 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>10.5,-25,15,-25</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12.5,-28.5,15,-28.5</points>
<connection>
<GID>40</GID>
<name>N_in0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>15,-27,20,-27</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>6,15.5,7,15.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,12,7,12</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-13.5,7,-9.5</points>
<intersection>-13.5 5</intersection>
<intersection>-9.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>7,-13.5,20.5,-13.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6,-9.5,7,-9.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>10.5,-15.5,20.5,-15.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>12.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12.5,-15.5,12.5,-12.5</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>-15.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-21.5,27.5,-10</points>
<intersection>-21.5 6</intersection>
<intersection>-14.5 1</intersection>
<intersection>-12 7</intersection>
<intersection>-10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-14.5,27.5,-14.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-10,27.5,-10</points>
<connection>
<GID>56</GID>
<name>N_in0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>27.5,-21.5,36.5,-21.5</points>
<connection>
<GID>70</GID>
<name>IN_B_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27.5,-12,33.5,-12</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-31,7,-29</points>
<intersection>-31 6</intersection>
<intersection>-29 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>7,-29,20,-29</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6,-31,7,-31</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-30,29,-21.5</points>
<intersection>-30 4</intersection>
<intersection>-28 5</intersection>
<intersection>-21.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26,-30,29,-30</points>
<intersection>26 7</intersection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>26,-28,29,-28</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>26,-31,26,-30</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<intersection>-30 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>29,-21.5,38.5,-21.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection>
<intersection>33.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>33.5,-21.5,33.5,-14</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>-21.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,-55,3.5,-54</points>
<intersection>-55 1</intersection>
<intersection>-54 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-55,4.5,-55</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-54,3.5,-54</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-31,37.5,-27.5</points>
<connection>
<GID>72</GID>
<name>N_in3</name></connection>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>-29 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>37.5,-29,49,-29</points>
<intersection>37.5 0</intersection>
<intersection>49 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>49,-29,49,-26</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>-29 5</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,15.5,20.5,15.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<connection>
<GID>74</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-0.5,-58,-0.5,-57</points>
<intersection>-58 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-0.5,-57,4.5,-57</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>-0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-58,-0.5,-58</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-59.5,15,-56</points>
<intersection>-59.5 9</intersection>
<intersection>-58 10</intersection>
<intersection>-56 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>10.5,-56,15,-56</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12.5,-59.5,15,-59.5</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>15,-58,20,-58</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-44.5,7,-40.5</points>
<intersection>-44.5 5</intersection>
<intersection>-40.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>7,-44.5,20.5,-44.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6,-40.5,7,-40.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-30,56.5,-18</points>
<intersection>-30 5</intersection>
<intersection>-25 6</intersection>
<intersection>-18 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56.5,-18,58.5,-18</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>55,-30,56.5,-30</points>
<connection>
<GID>90</GID>
<name>N_in0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>55,-25,56.5,-25</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,15.5,33,15.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>10.5,-46.5,20.5,-46.5</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>12.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12.5,-46.5,12.5,-43.5</points>
<connection>
<GID>9</GID>
<name>N_in0</name></connection>
<intersection>-46.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-52.5,27.5,-41</points>
<intersection>-52.5 6</intersection>
<intersection>-45.5 1</intersection>
<intersection>-43 7</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-45.5,27.5,-45.5</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-41,27.5,-41</points>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>27.5,-52.5,36.5,-52.5</points>
<connection>
<GID>33</GID>
<name>IN_B_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27.5,-43,33.5,-43</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-20.5,65.5,-17</points>
<connection>
<GID>104</GID>
<name>N_in3</name></connection>
<intersection>-18 3</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-17,65.5,-17</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>65.5,-18,69.5,-18</points>
<connection>
<GID>102</GID>
<name>IN_1</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-62,7,-60</points>
<intersection>-62 6</intersection>
<intersection>-60 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>7,-60,20,-60</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6,-62,7,-62</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-13,40,-7.5</points>
<intersection>-13 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-7.5,49,-7.5</points>
<connection>
<GID>68</GID>
<name>N_in0</name></connection>
<intersection>40 0</intersection>
<intersection>49 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-13,40,-13</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>40 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49,-9,49,-7.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-23.5,20.5,-20.5</points>
<intersection>-23.5 10</intersection>
<intersection>-20.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>20.5,-23.5,49,-23.5</points>
<intersection>20.5 0</intersection>
<intersection>41.5 12</intersection>
<intersection>49 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-8,-20.5,20.5,-20.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>41.5,-23.5,41.5,-17.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-23.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>49,-24,49,-23.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>-23.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-17.5,48,-11</points>
<intersection>-17.5 4</intersection>
<intersection>-11 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>48,-11,49,-11</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>47.5,-17.5,48,-17.5</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-16,56,-9</points>
<connection>
<GID>88</GID>
<name>N_in2</name></connection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-16,58.5,-16</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>55 3</intersection>
<intersection>56 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55,-16,55,-10</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>-16 1</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-61,29,-52.5</points>
<intersection>-61 4</intersection>
<intersection>-59 5</intersection>
<intersection>-52.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26,-61,29,-61</points>
<intersection>26 7</intersection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>26,-59,29,-59</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>26,-62,26,-61</points>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<intersection>-61 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>29,-52.5,38.5,-52.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection>
<intersection>33.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>33.5,-52.5,33.5,-45</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-52.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-16,31.5,-5.5</points>
<intersection>-16 12</intersection>
<intersection>-5.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>31.5,-16,69.5,-16</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-6,-5.5,31.5,-5.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81.5,-23.5,85,-23.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<connection>
<GID>116</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-23.5,91,-23.5</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<connection>
<GID>118</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-17,77.5,-17</points>
<connection>
<GID>102</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>N_in0</name></connection>
<intersection>75.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75.5,-27,75.5,-17</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>-27 3</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75.5,-27,76,-27</points>
<connection>
<GID>114</GID>
<name>N_in3</name></connection>
<intersection>75.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-62,37.5,-58.5</points>
<connection>
<GID>35</GID>
<name>N_in3</name></connection>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>-61 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>37.5,-61,49,-61</points>
<intersection>37.5 0</intersection>
<intersection>49 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>49,-61,49,-57</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-61 5</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-61,56.5,-49</points>
<intersection>-61 5</intersection>
<intersection>-56 6</intersection>
<intersection>-49 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56.5,-49,58.5,-49</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>55,-61,56.5,-61</points>
<connection>
<GID>49</GID>
<name>N_in0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>55,-56,56.5,-56</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-51.5,65.5,-48</points>
<connection>
<GID>54</GID>
<name>N_in3</name></connection>
<intersection>-49 3</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-48,65.5,-48</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>65.5,-49,69.5,-49</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-44,40,-38.5</points>
<intersection>-44 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-38.5,49,-38.5</points>
<connection>
<GID>31</GID>
<name>N_in0</name></connection>
<intersection>40 0</intersection>
<intersection>49 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-44,40,-44</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>40 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>49,-40,49,-38.5</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>-38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-54.5,20.5,-51.5</points>
<intersection>-54.5 10</intersection>
<intersection>-51.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>20.5,-54.5,49,-54.5</points>
<intersection>20.5 0</intersection>
<intersection>41.5 12</intersection>
<intersection>49 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-8,-51.5,20.5,-51.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>41.5,-54.5,41.5,-48.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-54.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>49,-55,49,-54.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-54.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-48.5,48,-42</points>
<intersection>-48.5 4</intersection>
<intersection>-42 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>48,-42,49,-42</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>47.5,-48.5,48,-48.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-47,56,-40</points>
<connection>
<GID>47</GID>
<name>N_in2</name></connection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-47,58.5,-47</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>55 3</intersection>
<intersection>56 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55,-47,55,-41</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>-47 1</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-47,31.5,-36.5</points>
<intersection>-47 12</intersection>
<intersection>-36.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>31.5,-47,69.5,-47</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-6,-36.5,31.5,-36.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81.5,-54.5,85,-54.5</points>
<connection>
<GID>57</GID>
<name>OUT</name></connection>
<connection>
<GID>61</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-54.5,91,-54.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<connection>
<GID>62</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-48,77.5,-48</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>55</GID>
<name>N_in0</name></connection>
<intersection>75.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75.5,-58,75.5,-48</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>-58 3</intersection>
<intersection>-48 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75.5,-58,76,-58</points>
<connection>
<GID>59</GID>
<name>N_in3</name></connection>
<intersection>75.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-74.5,-5,-74.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-75.5,2,-74.5</points>
<intersection>-75.5 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-75.5,4,-75.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-74.5,2,-74.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-78.5,-3.5,-77.5</points>
<intersection>-78.5 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,-77.5,4,-77.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-78.5,-3.5,-78.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-84,-4,-84</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<connection>
<GID>73</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-85,3,-84</points>
<intersection>-85 1</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-85,4,-85</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-84,3,-84</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-88,-1,-87</points>
<intersection>-88 2</intersection>
<intersection>-87 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-87,4,-87</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-88,-1,-88</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-89.5,14.5,-86</points>
<intersection>-89.5 9</intersection>
<intersection>-88 10</intersection>
<intersection>-86 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>10,-86,14.5,-86</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12,-89.5,14.5,-89.5</points>
<connection>
<GID>81</GID>
<name>N_in0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>14.5,-88,19.5,-88</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-74.5,6.5,-70.5</points>
<intersection>-74.5 5</intersection>
<intersection>-70.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-74.5,20,-74.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6.5,-70.5,6.5,-70.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>10,-76.5,20,-76.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>12 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12,-76.5,12,-73.5</points>
<connection>
<GID>71</GID>
<name>N_in0</name></connection>
<intersection>-76.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-82.5,27,-71</points>
<intersection>-82.5 6</intersection>
<intersection>-75.5 1</intersection>
<intersection>-73 7</intersection>
<intersection>-71 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-75.5,27,-75.5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-71,27,-71</points>
<connection>
<GID>87</GID>
<name>N_in0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>27,-82.5,36,-82.5</points>
<connection>
<GID>97</GID>
<name>IN_B_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27,-73,33,-73</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-92,6.5,-90</points>
<intersection>-92 6</intersection>
<intersection>-90 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-90,19.5,-90</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6.5,-92,6.5,-92</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-91,28.5,-82.5</points>
<intersection>-91 4</intersection>
<intersection>-89 5</intersection>
<intersection>-82.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25.5,-91,28.5,-91</points>
<intersection>25.5 7</intersection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>25.5,-89,28.5,-89</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25.5,-92,25.5,-91</points>
<connection>
<GID>93</GID>
<name>N_in0</name></connection>
<intersection>-91 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>28.5,-82.5,38,-82.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection>
<intersection>33 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>33,-82.5,33,-75</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>-82.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-92,37,-88.5</points>
<connection>
<GID>98</GID>
<name>N_in3</name></connection>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>-90.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>37,-90.5,48.5,-90.5</points>
<intersection>37 0</intersection>
<intersection>48.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>48.5,-90.5,48.5,-87</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>-90.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-91,56,-79</points>
<intersection>-91 5</intersection>
<intersection>-86 6</intersection>
<intersection>-79 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56,-79,58,-79</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54.5,-91,56,-91</points>
<connection>
<GID>108</GID>
<name>N_in0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54.5,-86,56,-86</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-81.5,65,-78</points>
<connection>
<GID>113</GID>
<name>N_in3</name></connection>
<intersection>-79 3</intersection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64,-78,65,-78</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>65 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>65,-79,69,-79</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-74,39.5,-68.5</points>
<intersection>-74 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-68.5,48.5,-68.5</points>
<connection>
<GID>96</GID>
<name>N_in0</name></connection>
<intersection>39.5 0</intersection>
<intersection>48.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-74,39.5,-74</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48.5,-70,48.5,-68.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>-68.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-84.5,20,-81.5</points>
<intersection>-84.5 10</intersection>
<intersection>-81.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>20,-84.5,48.5,-84.5</points>
<intersection>20 0</intersection>
<intersection>41 12</intersection>
<intersection>48.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-8.5,-81.5,20,-81.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>41,-84.5,41,-78.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-84.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>48.5,-85,48.5,-84.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-84.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-78.5,47.5,-72</points>
<intersection>-78.5 4</intersection>
<intersection>-72 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47.5,-72,48.5,-72</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>47,-78.5,47.5,-78.5</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-77,55.5,-70</points>
<connection>
<GID>107</GID>
<name>N_in2</name></connection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-77,58,-77</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection>
<intersection>55.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-77,54.5,-71</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<intersection>-77 1</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-77,31,-66.5</points>
<intersection>-77 12</intersection>
<intersection>-66.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>31,-77,69,-77</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-6.5,-66.5,31,-66.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-84.5,84.5,-84.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<connection>
<GID>117</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-84.5,90.5,-84.5</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<connection>
<GID>121</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-78,77,-78</points>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-88,75,-78</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-88 3</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-88,75.5,-88</points>
<connection>
<GID>119</GID>
<name>N_in3</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-104,-5,-104</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-105,2,-104</points>
<intersection>-105 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-105,4,-105</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-104,2,-104</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-108,-3.5,-107</points>
<intersection>-108 2</intersection>
<intersection>-107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,-107,4,-107</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-108,-3.5,-108</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-113.5,-4,-113.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-114.5,3,-113.5</points>
<intersection>-114.5 1</intersection>
<intersection>-113.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-114.5,4,-114.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-113.5,3,-113.5</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-117.5,-1,-116.5</points>
<intersection>-117.5 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-116.5,4,-116.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-117.5,-1,-117.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-119,14.5,-115.5</points>
<intersection>-119 9</intersection>
<intersection>-117.5 10</intersection>
<intersection>-115.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>10,-115.5,14.5,-115.5</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12,-119,14.5,-119</points>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>14.5,-117.5,19.5,-117.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-104,6.5,-100</points>
<intersection>-104 5</intersection>
<intersection>-100 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-104,20,-104</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6.5,-100,6.5,-100</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>10,-106,20,-106</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>12 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12,-106,12,-103</points>
<connection>
<GID>126</GID>
<name>N_in0</name></connection>
<intersection>-106 2</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-112,27,-100.5</points>
<intersection>-112 6</intersection>
<intersection>-105 1</intersection>
<intersection>-102.5 7</intersection>
<intersection>-100.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-105,27,-105</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-100.5,27,-100.5</points>
<connection>
<GID>134</GID>
<name>N_in0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>27,-112,36,-112</points>
<connection>
<GID>140</GID>
<name>IN_B_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27,-102.5,33,-102.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-121.5,6.5,-119.5</points>
<intersection>-121.5 6</intersection>
<intersection>-119.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-119.5,19.5,-119.5</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6.5,-121.5,6.5,-121.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-120.5,28.5,-112</points>
<intersection>-120.5 4</intersection>
<intersection>-118.5 5</intersection>
<intersection>-112 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25.5,-120.5,28.5,-120.5</points>
<intersection>25.5 7</intersection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>25.5,-118.5,28.5,-118.5</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25.5,-121.5,25.5,-120.5</points>
<connection>
<GID>137</GID>
<name>N_in0</name></connection>
<intersection>-120.5 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>28.5,-112,38,-112</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection>
<intersection>33 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>33,-112,33,-104.5</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-112 9</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-121.5,37,-118</points>
<connection>
<GID>141</GID>
<name>N_in3</name></connection>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>-121 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>37,-121,48.5,-121</points>
<intersection>37 0</intersection>
<intersection>48.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>48.5,-121,48.5,-116.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>-121 5</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-120.5,56,-108.5</points>
<intersection>-120.5 5</intersection>
<intersection>-115.5 6</intersection>
<intersection>-108.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56,-108.5,58,-108.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54.5,-120.5,56,-120.5</points>
<connection>
<GID>148</GID>
<name>N_in0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54.5,-115.5,56,-115.5</points>
<connection>
<GID>145</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-111,65,-107.5</points>
<connection>
<GID>151</GID>
<name>N_in3</name></connection>
<intersection>-108.5 3</intersection>
<intersection>-107.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64,-107.5,65,-107.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>65 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>65,-108.5,69,-108.5</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-103.5,39.5,-98</points>
<intersection>-103.5 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-98,48.5,-98</points>
<connection>
<GID>139</GID>
<name>N_in0</name></connection>
<intersection>39.5 0</intersection>
<intersection>48.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-103.5,39.5,-103.5</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48.5,-99.5,48.5,-98</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-98 1</intersection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-114,20,-111</points>
<intersection>-114 10</intersection>
<intersection>-111 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>20,-114,48.5,-114</points>
<intersection>20 0</intersection>
<intersection>41 12</intersection>
<intersection>48.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-8.5,-111,20,-111</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>41,-114,41,-108</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>-114 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>48.5,-114.5,48.5,-114</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-114 10</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-108,47.5,-101.5</points>
<intersection>-108 4</intersection>
<intersection>-101.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47.5,-101.5,48.5,-101.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>47,-108,47.5,-108</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-106.5,55.5,-99.5</points>
<connection>
<GID>147</GID>
<name>N_in2</name></connection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-106.5,58,-106.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection>
<intersection>55.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-106.5,54.5,-100.5</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>-106.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-106.5,31,-96</points>
<intersection>-106.5 12</intersection>
<intersection>-96 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>31,-106.5,69,-106.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-6.5,-96,31,-96</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-114,84.5,-114</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>153</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-114,90.5,-114</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<connection>
<GID>156</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-107.5,77,-107.5</points>
<connection>
<GID>152</GID>
<name>N_in0</name></connection>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-117.5,75,-107.5</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-117.5 3</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-117.5,75.5,-117.5</points>
<connection>
<GID>154</GID>
<name>N_in3</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-134,-5,-134</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<connection>
<GID>158</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-135,2,-134</points>
<intersection>-135 1</intersection>
<intersection>-134 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-135,4,-135</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-134,2,-134</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-138,-3.5,-137</points>
<intersection>-138 2</intersection>
<intersection>-137 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,-137,4,-137</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-138,-3.5,-138</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-143.5,-4,-143.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-144.5,3,-143.5</points>
<intersection>-144.5 1</intersection>
<intersection>-143.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-144.5,4,-144.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-143.5,3,-143.5</points>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-147.5,-1,-146.5</points>
<intersection>-147.5 2</intersection>
<intersection>-146.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-146.5,4,-146.5</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-147.5,-1,-147.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-149,14.5,-145.5</points>
<intersection>-149 9</intersection>
<intersection>-147.5 10</intersection>
<intersection>-145.5 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>10,-145.5,14.5,-145.5</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12,-149,14.5,-149</points>
<connection>
<GID>166</GID>
<name>N_in0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>14.5,-147.5,19.5,-147.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-134,6.5,-130</points>
<intersection>-134 5</intersection>
<intersection>-130 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-134,20,-134</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6.5,-130,6.5,-130</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>10,-136,20,-136</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>12 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12,-136,12,-133</points>
<connection>
<GID>161</GID>
<name>N_in0</name></connection>
<intersection>-136 2</intersection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-142,27,-130.5</points>
<intersection>-142 6</intersection>
<intersection>-135 1</intersection>
<intersection>-132.5 7</intersection>
<intersection>-130.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-135,27,-135</points>
<connection>
<GID>168</GID>
<name>OUT</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-130.5,27,-130.5</points>
<connection>
<GID>169</GID>
<name>N_in0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>27,-142,36,-142</points>
<connection>
<GID>175</GID>
<name>IN_B_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27,-132.5,33,-132.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-151.5,6.5,-149.5</points>
<intersection>-151.5 6</intersection>
<intersection>-149.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-149.5,19.5,-149.5</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6.5,-151.5,6.5,-151.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-150.5,28.5,-142</points>
<intersection>-150.5 4</intersection>
<intersection>-148.5 5</intersection>
<intersection>-142 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25.5,-150.5,28.5,-150.5</points>
<intersection>25.5 7</intersection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>25.5,-148.5,28.5,-148.5</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25.5,-151.5,25.5,-150.5</points>
<connection>
<GID>172</GID>
<name>N_in0</name></connection>
<intersection>-150.5 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>28.5,-142,38,-142</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection>
<intersection>33 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>33,-142,33,-134.5</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>-142 9</intersection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-151.5,37,-148</points>
<connection>
<GID>176</GID>
<name>N_in3</name></connection>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection>
<intersection>-150 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>37,-150,48.5,-150</points>
<intersection>37 0</intersection>
<intersection>48.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>48.5,-150,48.5,-146.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>-150 5</intersection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-150.5,56,-138.5</points>
<intersection>-150.5 5</intersection>
<intersection>-145.5 6</intersection>
<intersection>-138.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56,-138.5,58,-138.5</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54.5,-150.5,56,-150.5</points>
<connection>
<GID>183</GID>
<name>N_in0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54.5,-145.5,56,-145.5</points>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-141,65,-137.5</points>
<connection>
<GID>186</GID>
<name>N_in3</name></connection>
<intersection>-138.5 3</intersection>
<intersection>-137.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64,-137.5,65,-137.5</points>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<intersection>65 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>65,-138.5,69,-138.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-133.5,39.5,-128</points>
<intersection>-133.5 2</intersection>
<intersection>-128 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-128,48.5,-128</points>
<connection>
<GID>174</GID>
<name>N_in0</name></connection>
<intersection>39.5 0</intersection>
<intersection>48.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-133.5,39.5,-133.5</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48.5,-129.5,48.5,-128</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>-128 1</intersection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-144,20,-141</points>
<intersection>-144 10</intersection>
<intersection>-141 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>20,-144,48.5,-144</points>
<intersection>20 0</intersection>
<intersection>41 12</intersection>
<intersection>48.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-8.5,-141,20,-141</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>41,-144,41,-138</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>-144 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>48.5,-144.5,48.5,-144</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-144 10</intersection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-138,47.5,-131.5</points>
<intersection>-138 4</intersection>
<intersection>-131.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47.5,-131.5,48.5,-131.5</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>47,-138,47.5,-138</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-136.5,55.5,-129.5</points>
<connection>
<GID>182</GID>
<name>N_in2</name></connection>
<intersection>-136.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-136.5,58,-136.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection>
<intersection>55.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-136.5,54.5,-130.5</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>-136.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-136.5,31,-126</points>
<intersection>-136.5 12</intersection>
<intersection>-126 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>31,-136.5,69,-136.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-6.5,-126,31,-126</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-144,84.5,-144</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<connection>
<GID>188</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-144,90.5,-144</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<connection>
<GID>191</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-137.5,77,-137.5</points>
<connection>
<GID>187</GID>
<name>N_in0</name></connection>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-147.5,75,-137.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-147.5 3</intersection>
<intersection>-137.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-147.5,75.5,-147.5</points>
<connection>
<GID>189</GID>
<name>N_in3</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-163.5,-5,-163.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<connection>
<GID>193</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-164.5,2,-163.5</points>
<intersection>-164.5 1</intersection>
<intersection>-163.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-164.5,4,-164.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,-163.5,2,-163.5</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-167.5,-3.5,-166.5</points>
<intersection>-167.5 2</intersection>
<intersection>-166.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,-166.5,4,-166.5</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-167.5,-3.5,-167.5</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-6.5,-173,-4,-173</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<connection>
<GID>197</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-174,3,-173</points>
<intersection>-174 1</intersection>
<intersection>-173 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-174,4,-174</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2,-173,3,-173</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1,-177,-1,-176</points>
<intersection>-177 2</intersection>
<intersection>-176 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1,-176,4,-176</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>-1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-177,-1,-177</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>-1 0</intersection></hsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-178.5,14.5,-175</points>
<intersection>-178.5 9</intersection>
<intersection>-177 10</intersection>
<intersection>-175 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>10,-175,14.5,-175</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>12,-178.5,14.5,-178.5</points>
<connection>
<GID>201</GID>
<name>N_in0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>14.5,-177,19.5,-177</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-163.5,6.5,-159.5</points>
<intersection>-163.5 5</intersection>
<intersection>-159.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-163.5,20,-163.5</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6.5,-159.5,6.5,-159.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>10,-165.5,20,-165.5</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<intersection>12 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>12,-165.5,12,-162.5</points>
<connection>
<GID>196</GID>
<name>N_in0</name></connection>
<intersection>-165.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-171.5,27,-160</points>
<intersection>-171.5 6</intersection>
<intersection>-164.5 1</intersection>
<intersection>-162 7</intersection>
<intersection>-160 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-164.5,27,-164.5</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-160,27,-160</points>
<connection>
<GID>204</GID>
<name>N_in0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>27,-171.5,36,-171.5</points>
<connection>
<GID>210</GID>
<name>IN_B_0</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>27,-162,33,-162</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-181,6.5,-179</points>
<intersection>-181 6</intersection>
<intersection>-179 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>6.5,-179,19.5,-179</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-6.5,-181,6.5,-181</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-180,28.5,-171.5</points>
<intersection>-180 4</intersection>
<intersection>-178 5</intersection>
<intersection>-171.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>25.5,-180,28.5,-180</points>
<intersection>25.5 7</intersection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>25.5,-178,28.5,-178</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25.5,-181,25.5,-180</points>
<connection>
<GID>207</GID>
<name>N_in0</name></connection>
<intersection>-180 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>28.5,-171.5,38,-171.5</points>
<connection>
<GID>210</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection>
<intersection>33 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>33,-171.5,33,-164</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>-171.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-181,37,-177.5</points>
<connection>
<GID>211</GID>
<name>N_in3</name></connection>
<connection>
<GID>210</GID>
<name>OUT_0</name></connection>
<intersection>-180.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>37,-180.5,48.5,-180.5</points>
<intersection>37 0</intersection>
<intersection>48.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>48.5,-180.5,48.5,-176</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>-180.5 5</intersection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-180,56,-168</points>
<intersection>-180 5</intersection>
<intersection>-175 6</intersection>
<intersection>-168 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56,-168,58,-168</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54.5,-180,56,-180</points>
<connection>
<GID>218</GID>
<name>N_in0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>54.5,-175,56,-175</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-170.5,65,-167</points>
<connection>
<GID>221</GID>
<name>N_in3</name></connection>
<intersection>-168 3</intersection>
<intersection>-167 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>64,-167,65,-167</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<intersection>65 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>65,-168,69,-168</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-163,39.5,-157.5</points>
<intersection>-163 2</intersection>
<intersection>-157.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-157.5,48.5,-157.5</points>
<connection>
<GID>209</GID>
<name>N_in0</name></connection>
<intersection>39.5 0</intersection>
<intersection>48.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-163,39.5,-163</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48.5,-159,48.5,-157.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>-157.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-173.5,20,-170.5</points>
<intersection>-173.5 10</intersection>
<intersection>-170.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>20,-173.5,48.5,-173.5</points>
<intersection>20 0</intersection>
<intersection>41 12</intersection>
<intersection>48.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-8.5,-170.5,20,-170.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>41,-173.5,41,-167.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>-173.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>48.5,-174,48.5,-173.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>-173.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-167.5,47.5,-161</points>
<intersection>-167.5 4</intersection>
<intersection>-161 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>47.5,-161,48.5,-161</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>47.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>47,-167.5,47.5,-167.5</points>
<connection>
<GID>213</GID>
<name>OUT_0</name></connection>
<intersection>47.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-166,55.5,-159</points>
<connection>
<GID>217</GID>
<name>N_in2</name></connection>
<intersection>-166 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-166,58,-166</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection>
<intersection>55.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-166,54.5,-160</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>-166 1</intersection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-166,31,-155.5</points>
<intersection>-166 12</intersection>
<intersection>-155.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>31,-166,69,-166</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-6.5,-155.5,31,-155.5</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81,-173.5,84.5,-173.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<connection>
<GID>223</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-173.5,90.5,-173.5</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<connection>
<GID>226</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-167,77,-167</points>
<connection>
<GID>222</GID>
<name>N_in0</name></connection>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<intersection>75 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>75,-177,75,-167</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>-177 3</intersection>
<intersection>-167 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>75,-177,75.5,-177</points>
<connection>
<GID>224</GID>
<name>N_in3</name></connection>
<intersection>75 2</intersection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8.5,-196.5,-7,-196.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<connection>
<GID>229</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-197.5,0,-196.5</points>
<intersection>-197.5 1</intersection>
<intersection>-196.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0,-197.5,2,-197.5</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1,-196.5,0,-196.5</points>
<connection>
<GID>229</GID>
<name>OUT_0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-200.5,-5.5,-199.5</points>
<intersection>-200.5 2</intersection>
<intersection>-199.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-5.5,-199.5,2,-199.5</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<intersection>-5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,-200.5,-5.5,-200.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8.5,-206,-6,-206</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<connection>
<GID>234</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,-207,1,-206</points>
<intersection>-207 1</intersection>
<intersection>-206 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-207,2,-207</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-206,1,-206</points>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3,-210,-3,-209</points>
<intersection>-210 2</intersection>
<intersection>-209 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3,-209,2,-209</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<intersection>-3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-10,-210,-3,-210</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>-3 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-211.5,12.5,-208</points>
<intersection>-211.5 9</intersection>
<intersection>-210 10</intersection>
<intersection>-208 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>8,-208,12.5,-208</points>
<connection>
<GID>235</GID>
<name>OUT</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>10,-211.5,12.5,-211.5</points>
<connection>
<GID>236</GID>
<name>N_in0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>12.5,-210,17.5,-210</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-196.5,4.5,-192.5</points>
<intersection>-196.5 5</intersection>
<intersection>-192.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4.5,-196.5,18,-196.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-8.5,-192.5,4.5,-192.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>8,-198.5,18,-198.5</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>10 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>10,-198.5,10,-195.5</points>
<connection>
<GID>231</GID>
<name>N_in0</name></connection>
<intersection>-198.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-204.5,25,-193</points>
<intersection>-204.5 6</intersection>
<intersection>-197.5 1</intersection>
<intersection>-195 7</intersection>
<intersection>-193 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-197.5,25,-197.5</points>
<connection>
<GID>238</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-193,25,-193</points>
<connection>
<GID>239</GID>
<name>N_in0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>25,-204.5,34,-204.5</points>
<connection>
<GID>245</GID>
<name>IN_B_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>25,-195,31,-195</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>4.5,-214,4.5,-212</points>
<intersection>-214 6</intersection>
<intersection>-212 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>4.5,-212,17.5,-212</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<intersection>4.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-8.5,-214,4.5,-214</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-213,26.5,-204.5</points>
<intersection>-213 4</intersection>
<intersection>-211 5</intersection>
<intersection>-204.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>23.5,-213,26.5,-213</points>
<intersection>23.5 7</intersection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>23.5,-211,26.5,-211</points>
<connection>
<GID>241</GID>
<name>OUT</name></connection>
<intersection>26.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>23.5,-214,23.5,-213</points>
<connection>
<GID>242</GID>
<name>N_in0</name></connection>
<intersection>-213 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>26.5,-204.5,36,-204.5</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection>
<intersection>31 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>31,-204.5,31,-197</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>-204.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-214,35,-210.5</points>
<connection>
<GID>246</GID>
<name>N_in3</name></connection>
<connection>
<GID>245</GID>
<name>OUT_0</name></connection>
<intersection>-212 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>35,-212,46.5,-212</points>
<intersection>35 0</intersection>
<intersection>46.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>46.5,-212,46.5,-209</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>-212 5</intersection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-213,54,-201</points>
<intersection>-213 5</intersection>
<intersection>-208 6</intersection>
<intersection>-201 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>54,-201,56,-201</points>
<connection>
<GID>251</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>52.5,-213,54,-213</points>
<connection>
<GID>253</GID>
<name>N_in0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>52.5,-208,54,-208</points>
<connection>
<GID>250</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-203.5,63,-200</points>
<connection>
<GID>256</GID>
<name>N_in3</name></connection>
<intersection>-201 3</intersection>
<intersection>-200 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62,-200,63,-200</points>
<connection>
<GID>251</GID>
<name>OUT</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>63,-201,67,-201</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-196,37.5,-190.5</points>
<intersection>-196 2</intersection>
<intersection>-190.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-190.5,46.5,-190.5</points>
<connection>
<GID>244</GID>
<name>N_in0</name></connection>
<intersection>37.5 0</intersection>
<intersection>46.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-196,37.5,-196</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>46.5,-192,46.5,-190.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>-190.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-206.5,18,-203.5</points>
<intersection>-206.5 10</intersection>
<intersection>-203.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>18,-206.5,46.5,-206.5</points>
<intersection>18 0</intersection>
<intersection>39 12</intersection>
<intersection>46.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-10.5,-203.5,18,-203.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>39,-206.5,39,-200.5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>-206.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>46.5,-207,46.5,-206.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>-206.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-200.5,45.5,-194</points>
<intersection>-200.5 4</intersection>
<intersection>-194 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>45.5,-194,46.5,-194</points>
<connection>
<GID>249</GID>
<name>IN_1</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>45,-200.5,45.5,-200.5</points>
<connection>
<GID>248</GID>
<name>OUT_0</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-199,53.5,-192</points>
<connection>
<GID>252</GID>
<name>N_in2</name></connection>
<intersection>-199 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-199,56,-199</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>52.5 3</intersection>
<intersection>53.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52.5,-199,52.5,-193</points>
<connection>
<GID>249</GID>
<name>OUT</name></connection>
<intersection>-199 1</intersection></vsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-199,29,-188.5</points>
<intersection>-199 12</intersection>
<intersection>-188.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>29,-199,67,-199</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>-8.5,-188.5,29,-188.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79,-206.5,82.5,-206.5</points>
<connection>
<GID>258</GID>
<name>OUT</name></connection>
<connection>
<GID>260</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-206.5,88.5,-206.5</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<connection>
<GID>261</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73,-200,75,-200</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<connection>
<GID>257</GID>
<name>N_in0</name></connection>
<intersection>73 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>73,-210,73,-200</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>-210 3</intersection>
<intersection>-200 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>73,-210,73.5,-210</points>
<connection>
<GID>259</GID>
<name>N_in3</name></connection>
<intersection>73 2</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-15.5,135,-15.5</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<connection>
<GID>264</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>171</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-16.5,142,-15.5</points>
<intersection>-16.5 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-16.5,144,-16.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-15.5,142,-15.5</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>172</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-19.5,136.5,-18.5</points>
<intersection>-19.5 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,-18.5,144,-18.5</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-19.5,136.5,-19.5</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>173</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-25,136,-25</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<connection>
<GID>269</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>174</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-26,143,-25</points>
<intersection>-26 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-26,144,-26</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>142,-25,143,-25</points>
<connection>
<GID>269</GID>
<name>OUT_0</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>175</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-29,139,-28</points>
<intersection>-29 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,-28,144,-28</points>
<connection>
<GID>270</GID>
<name>IN_1</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-29,139,-29</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>176</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-30.5,154.5,-27</points>
<intersection>-30.5 9</intersection>
<intersection>-29 10</intersection>
<intersection>-27 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>150,-27,154.5,-27</points>
<connection>
<GID>270</GID>
<name>OUT</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>152,-30.5,154.5,-30.5</points>
<connection>
<GID>271</GID>
<name>N_in0</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>154.5,-29,159.5,-29</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>154.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-15.5,146.5,-11.5</points>
<intersection>-15.5 5</intersection>
<intersection>-11.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>146.5,-15.5,160,-15.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>133.5,-11.5,146.5,-11.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>178</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>150,-17.5,160,-17.5</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<intersection>152 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>152,-17.5,152,-14.5</points>
<connection>
<GID>266</GID>
<name>N_in0</name></connection>
<intersection>-17.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-23.5,167,-12</points>
<intersection>-23.5 6</intersection>
<intersection>-16.5 1</intersection>
<intersection>-14 7</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-16.5,167,-16.5</points>
<connection>
<GID>273</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166,-12,167,-12</points>
<connection>
<GID>274</GID>
<name>N_in0</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>167,-23.5,176,-23.5</points>
<connection>
<GID>280</GID>
<name>IN_B_0</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>167,-14,173,-14</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-33,146.5,-31</points>
<intersection>-33 6</intersection>
<intersection>-31 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>146.5,-31,159.5,-31</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>133.5,-33,146.5,-33</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-32,168.5,-23.5</points>
<intersection>-32 4</intersection>
<intersection>-30 5</intersection>
<intersection>-23.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>165.5,-32,168.5,-32</points>
<intersection>165.5 7</intersection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>165.5,-30,168.5,-30</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<intersection>168.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>165.5,-33,165.5,-32</points>
<connection>
<GID>277</GID>
<name>N_in0</name></connection>
<intersection>-32 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>168.5,-23.5,178,-23.5</points>
<connection>
<GID>280</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection>
<intersection>173 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>173,-23.5,173,-16</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>-23.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-33,177,-29.5</points>
<connection>
<GID>281</GID>
<name>N_in3</name></connection>
<connection>
<GID>280</GID>
<name>OUT_0</name></connection>
<intersection>-32 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>177,-32,188.5,-32</points>
<intersection>177 0</intersection>
<intersection>188.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>188.5,-32,188.5,-28</points>
<connection>
<GID>285</GID>
<name>IN_1</name></connection>
<intersection>-32 5</intersection></vsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196,-32,196,-20</points>
<intersection>-32 5</intersection>
<intersection>-27 6</intersection>
<intersection>-20 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>196,-20,198,-20</points>
<connection>
<GID>286</GID>
<name>IN_1</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>194.5,-32,196,-32</points>
<connection>
<GID>288</GID>
<name>N_in0</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>194.5,-27,196,-27</points>
<connection>
<GID>285</GID>
<name>OUT</name></connection>
<intersection>196 0</intersection></hsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,-22.5,205,-19</points>
<connection>
<GID>291</GID>
<name>N_in3</name></connection>
<intersection>-20 3</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>204,-19,205,-19</points>
<connection>
<GID>286</GID>
<name>OUT</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>205,-20,209,-20</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<intersection>205 0</intersection></hsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-15,179.5,-9.5</points>
<intersection>-15 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179.5,-9.5,188.5,-9.5</points>
<connection>
<GID>279</GID>
<name>N_in0</name></connection>
<intersection>179.5 0</intersection>
<intersection>188.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179,-15,179.5,-15</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>179.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>188.5,-11,188.5,-9.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>-9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-25.5,160,-22.5</points>
<intersection>-25.5 10</intersection>
<intersection>-22.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>160,-25.5,188.5,-25.5</points>
<intersection>160 0</intersection>
<intersection>181 12</intersection>
<intersection>188.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>131.5,-22.5,160,-22.5</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>181,-25.5,181,-19.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>-25.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>188.5,-26,188.5,-25.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>-25.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-19.5,187.5,-13</points>
<intersection>-19.5 4</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>187.5,-13,188.5,-13</points>
<connection>
<GID>284</GID>
<name>IN_1</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>187,-19.5,187.5,-19.5</points>
<connection>
<GID>283</GID>
<name>OUT_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-18,195.5,-11</points>
<connection>
<GID>287</GID>
<name>N_in2</name></connection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194.5,-18,198,-18</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>194.5 3</intersection>
<intersection>195.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>194.5,-18,194.5,-12</points>
<connection>
<GID>284</GID>
<name>OUT</name></connection>
<intersection>-18 1</intersection></vsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-18,171,-7.5</points>
<intersection>-18 12</intersection>
<intersection>-7.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>171,-18,209,-18</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<intersection>171 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>133.5,-7.5,171,-7.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,-25.5,224.5,-25.5</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<connection>
<GID>295</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-25.5,230.5,-25.5</points>
<connection>
<GID>295</GID>
<name>OUT_0</name></connection>
<connection>
<GID>296</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-19,217,-19</points>
<connection>
<GID>290</GID>
<name>OUT</name></connection>
<connection>
<GID>292</GID>
<name>N_in0</name></connection>
<intersection>215 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>215,-29,215,-19</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>-29 3</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215,-29,215.5,-29</points>
<connection>
<GID>294</GID>
<name>N_in3</name></connection>
<intersection>215 2</intersection></hsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-46.5,135,-46.5</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<connection>
<GID>298</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-47.5,142,-46.5</points>
<intersection>-47.5 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-47.5,144,-47.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-46.5,142,-46.5</points>
<connection>
<GID>299</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-50.5,136.5,-49.5</points>
<intersection>-50.5 2</intersection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,-49.5,144,-49.5</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-50.5,136.5,-50.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-56,136,-56</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<connection>
<GID>302</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-57,143,-56</points>
<intersection>-57 1</intersection>
<intersection>-56 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-57,144,-57</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>142,-56,143,-56</points>
<connection>
<GID>304</GID>
<name>OUT_0</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-60,139,-59</points>
<intersection>-60 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,-59,144,-59</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-60,139,-60</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-61.5,154.5,-58</points>
<intersection>-61.5 9</intersection>
<intersection>-60 10</intersection>
<intersection>-58 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>150,-58,154.5,-58</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>152,-61.5,154.5,-61.5</points>
<connection>
<GID>306</GID>
<name>N_in0</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>154.5,-60,159.5,-60</points>
<connection>
<GID>311</GID>
<name>IN_0</name></connection>
<intersection>154.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-46.5,146.5,-42.5</points>
<intersection>-46.5 5</intersection>
<intersection>-42.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>146.5,-46.5,160,-46.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>133.5,-42.5,146.5,-42.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>150,-48.5,160,-48.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<intersection>152 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>152,-48.5,152,-45.5</points>
<connection>
<GID>301</GID>
<name>N_in0</name></connection>
<intersection>-48.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-54.5,167,-43</points>
<intersection>-54.5 6</intersection>
<intersection>-47.5 1</intersection>
<intersection>-45 7</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-47.5,167,-47.5</points>
<connection>
<GID>308</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166,-43,167,-43</points>
<connection>
<GID>309</GID>
<name>N_in0</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>167,-54.5,176,-54.5</points>
<connection>
<GID>315</GID>
<name>IN_B_0</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>167,-45,173,-45</points>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-64,146.5,-62</points>
<intersection>-64 6</intersection>
<intersection>-62 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>146.5,-62,159.5,-62</points>
<connection>
<GID>311</GID>
<name>IN_1</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>133.5,-64,146.5,-64</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-63,168.5,-54.5</points>
<intersection>-63 4</intersection>
<intersection>-61 5</intersection>
<intersection>-54.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>165.5,-63,168.5,-63</points>
<intersection>165.5 7</intersection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>165.5,-61,168.5,-61</points>
<connection>
<GID>311</GID>
<name>OUT</name></connection>
<intersection>168.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>165.5,-64,165.5,-63</points>
<connection>
<GID>312</GID>
<name>N_in0</name></connection>
<intersection>-63 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>168.5,-54.5,178,-54.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection>
<intersection>173 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>173,-54.5,173,-47</points>
<connection>
<GID>313</GID>
<name>IN_1</name></connection>
<intersection>-54.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-64,177,-60.5</points>
<connection>
<GID>316</GID>
<name>N_in3</name></connection>
<connection>
<GID>315</GID>
<name>OUT_0</name></connection>
<intersection>-63 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>177,-63,188.5,-63</points>
<intersection>177 0</intersection>
<intersection>188.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>188.5,-63,188.5,-59</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<intersection>-63 5</intersection></vsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196,-63,196,-51</points>
<intersection>-63 5</intersection>
<intersection>-58 6</intersection>
<intersection>-51 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>196,-51,198,-51</points>
<connection>
<GID>321</GID>
<name>IN_1</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>194.5,-63,196,-63</points>
<connection>
<GID>323</GID>
<name>N_in0</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>194.5,-58,196,-58</points>
<connection>
<GID>320</GID>
<name>OUT</name></connection>
<intersection>196 0</intersection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,-53.5,205,-50</points>
<connection>
<GID>326</GID>
<name>N_in3</name></connection>
<intersection>-51 3</intersection>
<intersection>-50 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>204,-50,205,-50</points>
<connection>
<GID>321</GID>
<name>OUT</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>205,-51,209,-51</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<intersection>205 0</intersection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-46,179.5,-40.5</points>
<intersection>-46 2</intersection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179.5,-40.5,188.5,-40.5</points>
<connection>
<GID>314</GID>
<name>N_in0</name></connection>
<intersection>179.5 0</intersection>
<intersection>188.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179,-46,179.5,-46</points>
<connection>
<GID>313</GID>
<name>OUT</name></connection>
<intersection>179.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>188.5,-42,188.5,-40.5</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>-40.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-56.5,160,-53.5</points>
<intersection>-56.5 10</intersection>
<intersection>-53.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>160,-56.5,188.5,-56.5</points>
<intersection>160 0</intersection>
<intersection>181 12</intersection>
<intersection>188.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>131.5,-53.5,160,-53.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>181,-56.5,181,-50.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>-56.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>188.5,-57,188.5,-56.5</points>
<connection>
<GID>320</GID>
<name>IN_0</name></connection>
<intersection>-56.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-50.5,187.5,-44</points>
<intersection>-50.5 4</intersection>
<intersection>-44 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>187.5,-44,188.5,-44</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>187,-50.5,187.5,-50.5</points>
<connection>
<GID>318</GID>
<name>OUT_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-49,195.5,-42</points>
<connection>
<GID>322</GID>
<name>N_in2</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194.5,-49,198,-49</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>194.5 3</intersection>
<intersection>195.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>194.5,-49,194.5,-43</points>
<connection>
<GID>319</GID>
<name>OUT</name></connection>
<intersection>-49 1</intersection></vsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-49,171,-38.5</points>
<intersection>-49 12</intersection>
<intersection>-38.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>171,-49,209,-49</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>171 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>133.5,-38.5,171,-38.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>213</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,-56.5,224.5,-56.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<connection>
<GID>328</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>214</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-56.5,230.5,-56.5</points>
<connection>
<GID>330</GID>
<name>OUT_0</name></connection>
<connection>
<GID>331</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>215</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-50,217,-50</points>
<connection>
<GID>327</GID>
<name>N_in0</name></connection>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<intersection>215 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>215,-60,215,-50</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>-60 3</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215,-60,215.5,-60</points>
<connection>
<GID>329</GID>
<name>N_in3</name></connection>
<intersection>215 2</intersection></hsegment></shape></wire>
<wire>
<ID>216</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134.5,-78.5,136,-78.5</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<connection>
<GID>333</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>217</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-79.5,143,-78.5</points>
<intersection>-79.5 1</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-79.5,145,-79.5</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>142,-78.5,143,-78.5</points>
<connection>
<GID>334</GID>
<name>OUT_0</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-82.5,137.5,-81.5</points>
<intersection>-82.5 2</intersection>
<intersection>-81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,-81.5,145,-81.5</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<intersection>137.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133,-82.5,137.5,-82.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134.5,-88,137,-88</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<connection>
<GID>337</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-89,144,-88</points>
<intersection>-89 1</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-89,145,-89</points>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-88,144,-88</points>
<connection>
<GID>339</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140,-92,140,-91</points>
<intersection>-92 2</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>140,-91,145,-91</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>140 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>133,-92,140,-92</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>140 0</intersection></hsegment></shape></wire>
<wire>
<ID>222</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155.5,-93.5,155.5,-90</points>
<intersection>-93.5 9</intersection>
<intersection>-92 10</intersection>
<intersection>-90 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>151,-90,155.5,-90</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>153,-93.5,155.5,-93.5</points>
<connection>
<GID>341</GID>
<name>N_in0</name></connection>
<intersection>155.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>155.5,-92,160.5,-92</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>155.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>223</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-78.5,147.5,-74.5</points>
<intersection>-78.5 5</intersection>
<intersection>-74.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>147.5,-78.5,161,-78.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>134.5,-74.5,147.5,-74.5</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>151,-80.5,161,-80.5</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<connection>
<GID>335</GID>
<name>OUT</name></connection>
<intersection>153 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>153,-80.5,153,-77.5</points>
<connection>
<GID>336</GID>
<name>N_in0</name></connection>
<intersection>-80.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168,-86.5,168,-75</points>
<intersection>-86.5 6</intersection>
<intersection>-79.5 1</intersection>
<intersection>-77 7</intersection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>167,-79.5,168,-79.5</points>
<connection>
<GID>343</GID>
<name>OUT</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,-75,168,-75</points>
<connection>
<GID>344</GID>
<name>N_in0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>168,-86.5,177,-86.5</points>
<connection>
<GID>350</GID>
<name>IN_B_0</name></connection>
<intersection>168 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>168,-77,174,-77</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<intersection>168 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-96,147.5,-94</points>
<intersection>-96 6</intersection>
<intersection>-94 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>147.5,-94,160.5,-94</points>
<connection>
<GID>346</GID>
<name>IN_1</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>134.5,-96,147.5,-96</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169.5,-95,169.5,-86.5</points>
<intersection>-95 4</intersection>
<intersection>-93 5</intersection>
<intersection>-86.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>166.5,-95,169.5,-95</points>
<intersection>166.5 7</intersection>
<intersection>169.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>166.5,-93,169.5,-93</points>
<connection>
<GID>346</GID>
<name>OUT</name></connection>
<intersection>169.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>166.5,-96,166.5,-95</points>
<connection>
<GID>347</GID>
<name>N_in0</name></connection>
<intersection>-95 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>169.5,-86.5,179,-86.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>169.5 0</intersection>
<intersection>174 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>174,-86.5,174,-79</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<intersection>-86.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178,-96,178,-92.5</points>
<connection>
<GID>351</GID>
<name>N_in3</name></connection>
<connection>
<GID>350</GID>
<name>OUT_0</name></connection>
<intersection>-93 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>178,-93,189.5,-93</points>
<intersection>178 0</intersection>
<intersection>189.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>189.5,-93,189.5,-91</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<intersection>-93 5</intersection></vsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197,-95,197,-83</points>
<intersection>-95 5</intersection>
<intersection>-90 6</intersection>
<intersection>-83 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>197,-83,199,-83</points>
<connection>
<GID>356</GID>
<name>IN_1</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>195.5,-95,197,-95</points>
<connection>
<GID>358</GID>
<name>N_in0</name></connection>
<intersection>197 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>195.5,-90,197,-90</points>
<connection>
<GID>355</GID>
<name>OUT</name></connection>
<intersection>197 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206,-85.5,206,-82</points>
<connection>
<GID>361</GID>
<name>N_in3</name></connection>
<intersection>-83 3</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>205,-82,206,-82</points>
<connection>
<GID>356</GID>
<name>OUT</name></connection>
<intersection>206 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>206,-83,210,-83</points>
<connection>
<GID>360</GID>
<name>IN_1</name></connection>
<intersection>206 0</intersection></hsegment></shape></wire>
<wire>
<ID>231</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>180.5,-78,180.5,-72.5</points>
<intersection>-78 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>180.5,-72.5,189.5,-72.5</points>
<connection>
<GID>349</GID>
<name>N_in0</name></connection>
<intersection>180.5 0</intersection>
<intersection>189.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>180,-78,180.5,-78</points>
<connection>
<GID>348</GID>
<name>OUT</name></connection>
<intersection>180.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>189.5,-74,189.5,-72.5</points>
<connection>
<GID>354</GID>
<name>IN_0</name></connection>
<intersection>-72.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>232</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-88.5,161,-85.5</points>
<intersection>-88.5 10</intersection>
<intersection>-85.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>161,-88.5,189.5,-88.5</points>
<intersection>161 0</intersection>
<intersection>182 12</intersection>
<intersection>189.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>132.5,-85.5,161,-85.5</points>
<connection>
<GID>352</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>182,-88.5,182,-82.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>-88.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>189.5,-89,189.5,-88.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>-88.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>233</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-82.5,188.5,-76</points>
<intersection>-82.5 4</intersection>
<intersection>-76 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>188.5,-76,189.5,-76</points>
<connection>
<GID>354</GID>
<name>IN_1</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>188,-82.5,188.5,-82.5</points>
<connection>
<GID>353</GID>
<name>OUT_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>234</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,-81,196.5,-74</points>
<connection>
<GID>357</GID>
<name>N_in2</name></connection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,-81,199,-81</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>195.5 3</intersection>
<intersection>196.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>195.5,-81,195.5,-75</points>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<intersection>-81 1</intersection></vsegment></shape></wire>
<wire>
<ID>235</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>172,-81,172,-70.5</points>
<intersection>-81 12</intersection>
<intersection>-70.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>172,-81,210,-81</points>
<connection>
<GID>360</GID>
<name>IN_0</name></connection>
<intersection>172 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>134.5,-70.5,172,-70.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>172 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>222,-88.5,225.5,-88.5</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<connection>
<GID>363</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>231.5,-88.5,231.5,-88.5</points>
<connection>
<GID>365</GID>
<name>OUT_0</name></connection>
<connection>
<GID>366</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>238</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>216,-82,218,-82</points>
<connection>
<GID>362</GID>
<name>N_in0</name></connection>
<connection>
<GID>360</GID>
<name>OUT</name></connection>
<intersection>216 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>216,-92,216,-82</points>
<connection>
<GID>363</GID>
<name>IN_1</name></connection>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<intersection>-92 3</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>216,-92,216.5,-92</points>
<connection>
<GID>364</GID>
<name>N_in3</name></connection>
<intersection>216 2</intersection></hsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135.5,-109.5,137,-109.5</points>
<connection>
<GID>369</GID>
<name>IN_0</name></connection>
<connection>
<GID>368</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-110.5,144,-109.5</points>
<intersection>-110.5 1</intersection>
<intersection>-109.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-110.5,146,-110.5</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-109.5,144,-109.5</points>
<connection>
<GID>369</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-113.5,138.5,-112.5</points>
<intersection>-113.5 2</intersection>
<intersection>-112.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-112.5,146,-112.5</points>
<connection>
<GID>370</GID>
<name>IN_1</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134,-113.5,138.5,-113.5</points>
<connection>
<GID>367</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135.5,-119,138,-119</points>
<connection>
<GID>374</GID>
<name>IN_0</name></connection>
<connection>
<GID>372</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-120,145,-119</points>
<intersection>-120 1</intersection>
<intersection>-119 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-120,146,-120</points>
<connection>
<GID>375</GID>
<name>IN_0</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144,-119,145,-119</points>
<connection>
<GID>374</GID>
<name>OUT_0</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-123,141,-122</points>
<intersection>-123 2</intersection>
<intersection>-122 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-122,146,-122</points>
<connection>
<GID>375</GID>
<name>IN_1</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134,-123,141,-123</points>
<connection>
<GID>373</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-124.5,156.5,-121</points>
<intersection>-124.5 9</intersection>
<intersection>-123 10</intersection>
<intersection>-121 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>152,-121,156.5,-121</points>
<connection>
<GID>375</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>154,-124.5,156.5,-124.5</points>
<connection>
<GID>376</GID>
<name>N_in0</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>156.5,-123,161.5,-123</points>
<connection>
<GID>381</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-109.5,148.5,-105.5</points>
<intersection>-109.5 5</intersection>
<intersection>-105.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>148.5,-109.5,162,-109.5</points>
<connection>
<GID>378</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>135.5,-105.5,148.5,-105.5</points>
<connection>
<GID>377</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>152,-111.5,162,-111.5</points>
<connection>
<GID>378</GID>
<name>IN_1</name></connection>
<connection>
<GID>370</GID>
<name>OUT</name></connection>
<intersection>154 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>154,-111.5,154,-108.5</points>
<connection>
<GID>371</GID>
<name>N_in0</name></connection>
<intersection>-111.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-117.5,169,-106</points>
<intersection>-117.5 6</intersection>
<intersection>-110.5 1</intersection>
<intersection>-108 7</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-110.5,169,-110.5</points>
<connection>
<GID>378</GID>
<name>OUT</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168,-106,169,-106</points>
<connection>
<GID>379</GID>
<name>N_in0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>169,-117.5,178,-117.5</points>
<connection>
<GID>385</GID>
<name>IN_B_0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>169,-108,175,-108</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-127,148.5,-125</points>
<intersection>-127 6</intersection>
<intersection>-125 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>148.5,-125,161.5,-125</points>
<connection>
<GID>381</GID>
<name>IN_1</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>135.5,-127,148.5,-127</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-126,170.5,-117.5</points>
<intersection>-126 4</intersection>
<intersection>-124 5</intersection>
<intersection>-117.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>167.5,-126,170.5,-126</points>
<intersection>167.5 7</intersection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>167.5,-124,170.5,-124</points>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<intersection>170.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>167.5,-127,167.5,-126</points>
<connection>
<GID>382</GID>
<name>N_in0</name></connection>
<intersection>-126 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>170.5,-117.5,180,-117.5</points>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection>
<intersection>175 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>175,-117.5,175,-110</points>
<connection>
<GID>383</GID>
<name>IN_1</name></connection>
<intersection>-117.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-127,179,-123.5</points>
<connection>
<GID>386</GID>
<name>N_in3</name></connection>
<connection>
<GID>385</GID>
<name>OUT_0</name></connection>
<intersection>-126 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>179,-126,190.5,-126</points>
<intersection>179 0</intersection>
<intersection>190.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>190.5,-126,190.5,-122</points>
<connection>
<GID>390</GID>
<name>IN_1</name></connection>
<intersection>-126 5</intersection></vsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-126,198,-114</points>
<intersection>-126 5</intersection>
<intersection>-121 6</intersection>
<intersection>-114 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>198,-114,200,-114</points>
<connection>
<GID>391</GID>
<name>IN_1</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>196.5,-126,198,-126</points>
<connection>
<GID>393</GID>
<name>N_in0</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>196.5,-121,198,-121</points>
<connection>
<GID>390</GID>
<name>OUT</name></connection>
<intersection>198 0</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-116.5,207,-113</points>
<connection>
<GID>396</GID>
<name>N_in3</name></connection>
<intersection>-114 3</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>206,-113,207,-113</points>
<connection>
<GID>391</GID>
<name>OUT</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207,-114,211,-114</points>
<connection>
<GID>395</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-109,181.5,-103.5</points>
<intersection>-109 2</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181.5,-103.5,190.5,-103.5</points>
<connection>
<GID>384</GID>
<name>N_in0</name></connection>
<intersection>181.5 0</intersection>
<intersection>190.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181,-109,181.5,-109</points>
<connection>
<GID>383</GID>
<name>OUT</name></connection>
<intersection>181.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>190.5,-105,190.5,-103.5</points>
<connection>
<GID>389</GID>
<name>IN_0</name></connection>
<intersection>-103.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-119.5,162,-116.5</points>
<intersection>-119.5 10</intersection>
<intersection>-116.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>162,-119.5,190.5,-119.5</points>
<intersection>162 0</intersection>
<intersection>183 12</intersection>
<intersection>190.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>133.5,-116.5,162,-116.5</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>183,-119.5,183,-113.5</points>
<connection>
<GID>388</GID>
<name>IN_0</name></connection>
<intersection>-119.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>190.5,-120,190.5,-119.5</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<intersection>-119.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,-113.5,189.5,-107</points>
<intersection>-113.5 4</intersection>
<intersection>-107 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189.5,-107,190.5,-107</points>
<connection>
<GID>389</GID>
<name>IN_1</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>189,-113.5,189.5,-113.5</points>
<connection>
<GID>388</GID>
<name>OUT_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-112,197.5,-105</points>
<connection>
<GID>392</GID>
<name>N_in2</name></connection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196.5,-112,200,-112</points>
<connection>
<GID>391</GID>
<name>IN_0</name></connection>
<intersection>196.5 3</intersection>
<intersection>197.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>196.5,-112,196.5,-106</points>
<connection>
<GID>389</GID>
<name>OUT</name></connection>
<intersection>-112 1</intersection></vsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-112,173,-101.5</points>
<intersection>-112 12</intersection>
<intersection>-101.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>173,-112,211,-112</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>135.5,-101.5,173,-101.5</points>
<connection>
<GID>394</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>223,-119.5,226.5,-119.5</points>
<connection>
<GID>400</GID>
<name>IN_0</name></connection>
<connection>
<GID>398</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-119.5,232.5,-119.5</points>
<connection>
<GID>400</GID>
<name>OUT_0</name></connection>
<connection>
<GID>401</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-113,219,-113</points>
<connection>
<GID>397</GID>
<name>N_in0</name></connection>
<connection>
<GID>395</GID>
<name>OUT</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-123,217,-113</points>
<connection>
<GID>398</GID>
<name>IN_1</name></connection>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<intersection>-123 3</intersection>
<intersection>-113 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-123,217.5,-123</points>
<connection>
<GID>399</GID>
<name>N_in3</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135.5,-140.5,137,-140.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<connection>
<GID>403</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144,-141.5,144,-140.5</points>
<intersection>-141.5 1</intersection>
<intersection>-140.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144,-141.5,146,-141.5</points>
<connection>
<GID>405</GID>
<name>IN_0</name></connection>
<intersection>144 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-140.5,144,-140.5</points>
<connection>
<GID>404</GID>
<name>OUT_0</name></connection>
<intersection>144 0</intersection></hsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-144.5,138.5,-143.5</points>
<intersection>-144.5 2</intersection>
<intersection>-143.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-143.5,146,-143.5</points>
<connection>
<GID>405</GID>
<name>IN_1</name></connection>
<intersection>138.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134,-144.5,138.5,-144.5</points>
<connection>
<GID>402</GID>
<name>IN_0</name></connection>
<intersection>138.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>135.5,-150,138,-150</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<connection>
<GID>407</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-151,145,-150</points>
<intersection>-151 1</intersection>
<intersection>-150 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-151,146,-151</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144,-150,145,-150</points>
<connection>
<GID>409</GID>
<name>OUT_0</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-154,141,-153</points>
<intersection>-154 2</intersection>
<intersection>-153 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-153,146,-153</points>
<connection>
<GID>410</GID>
<name>IN_1</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134,-154,141,-154</points>
<connection>
<GID>408</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-155.5,156.5,-152</points>
<intersection>-155.5 9</intersection>
<intersection>-154 10</intersection>
<intersection>-152 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>152,-152,156.5,-152</points>
<connection>
<GID>410</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>154,-155.5,156.5,-155.5</points>
<connection>
<GID>411</GID>
<name>N_in0</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>156.5,-154,161.5,-154</points>
<connection>
<GID>416</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-140.5,148.5,-136.5</points>
<intersection>-140.5 5</intersection>
<intersection>-136.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>148.5,-140.5,162,-140.5</points>
<connection>
<GID>413</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>135.5,-136.5,148.5,-136.5</points>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>152,-142.5,162,-142.5</points>
<connection>
<GID>413</GID>
<name>IN_1</name></connection>
<connection>
<GID>405</GID>
<name>OUT</name></connection>
<intersection>154 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>154,-142.5,154,-139.5</points>
<connection>
<GID>406</GID>
<name>N_in0</name></connection>
<intersection>-142.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>271</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>169,-148.5,169,-137</points>
<intersection>-148.5 6</intersection>
<intersection>-141.5 1</intersection>
<intersection>-139 7</intersection>
<intersection>-137 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>168,-141.5,169,-141.5</points>
<connection>
<GID>413</GID>
<name>OUT</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>168,-137,169,-137</points>
<connection>
<GID>414</GID>
<name>N_in0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>169,-148.5,178,-148.5</points>
<connection>
<GID>420</GID>
<name>IN_B_0</name></connection>
<intersection>169 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>169,-139,175,-139</points>
<connection>
<GID>418</GID>
<name>IN_0</name></connection>
<intersection>169 0</intersection></hsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148.5,-158,148.5,-156</points>
<intersection>-158 6</intersection>
<intersection>-156 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>148.5,-156,161.5,-156</points>
<connection>
<GID>416</GID>
<name>IN_1</name></connection>
<intersection>148.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>135.5,-158,148.5,-158</points>
<connection>
<GID>415</GID>
<name>IN_0</name></connection>
<intersection>148.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-157,170.5,-148.5</points>
<intersection>-157 4</intersection>
<intersection>-155 5</intersection>
<intersection>-148.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>167.5,-157,170.5,-157</points>
<intersection>167.5 7</intersection>
<intersection>170.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>167.5,-155,170.5,-155</points>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<intersection>170.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>167.5,-158,167.5,-157</points>
<connection>
<GID>417</GID>
<name>N_in0</name></connection>
<intersection>-157 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>170.5,-148.5,180,-148.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<intersection>170.5 0</intersection>
<intersection>175 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>175,-148.5,175,-141</points>
<connection>
<GID>418</GID>
<name>IN_1</name></connection>
<intersection>-148.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-158,179,-154.5</points>
<connection>
<GID>421</GID>
<name>N_in3</name></connection>
<connection>
<GID>420</GID>
<name>OUT_0</name></connection>
<intersection>-155 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>179,-155,190.5,-155</points>
<intersection>179 0</intersection>
<intersection>190.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>190.5,-155,190.5,-153</points>
<connection>
<GID>425</GID>
<name>IN_1</name></connection>
<intersection>-155 5</intersection></vsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-157,198,-145</points>
<intersection>-157 5</intersection>
<intersection>-152 6</intersection>
<intersection>-145 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>198,-145,200,-145</points>
<connection>
<GID>426</GID>
<name>IN_1</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>196.5,-157,198,-157</points>
<connection>
<GID>428</GID>
<name>N_in0</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>196.5,-152,198,-152</points>
<connection>
<GID>425</GID>
<name>OUT</name></connection>
<intersection>198 0</intersection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-147.5,207,-144</points>
<connection>
<GID>431</GID>
<name>N_in3</name></connection>
<intersection>-145 3</intersection>
<intersection>-144 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>206,-144,207,-144</points>
<connection>
<GID>426</GID>
<name>OUT</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>207,-145,211,-145</points>
<connection>
<GID>430</GID>
<name>IN_1</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>181.5,-140,181.5,-134.5</points>
<intersection>-140 2</intersection>
<intersection>-134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181.5,-134.5,190.5,-134.5</points>
<connection>
<GID>419</GID>
<name>N_in0</name></connection>
<intersection>181.5 0</intersection>
<intersection>190.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>181,-140,181.5,-140</points>
<connection>
<GID>418</GID>
<name>OUT</name></connection>
<intersection>181.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>190.5,-136,190.5,-134.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<intersection>-134.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>162,-150.5,162,-147.5</points>
<intersection>-150.5 10</intersection>
<intersection>-147.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>162,-150.5,190.5,-150.5</points>
<intersection>162 0</intersection>
<intersection>183 12</intersection>
<intersection>190.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>133.5,-147.5,162,-147.5</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<intersection>162 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>183,-150.5,183,-144.5</points>
<connection>
<GID>423</GID>
<name>IN_0</name></connection>
<intersection>-150.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>190.5,-151,190.5,-150.5</points>
<connection>
<GID>425</GID>
<name>IN_0</name></connection>
<intersection>-150.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189.5,-144.5,189.5,-138</points>
<intersection>-144.5 4</intersection>
<intersection>-138 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>189.5,-138,190.5,-138</points>
<connection>
<GID>424</GID>
<name>IN_1</name></connection>
<intersection>189.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>189,-144.5,189.5,-144.5</points>
<connection>
<GID>423</GID>
<name>OUT_0</name></connection>
<intersection>189.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>197.5,-143,197.5,-136</points>
<connection>
<GID>427</GID>
<name>N_in2</name></connection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196.5,-143,200,-143</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<intersection>196.5 3</intersection>
<intersection>197.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>196.5,-143,196.5,-137</points>
<connection>
<GID>424</GID>
<name>OUT</name></connection>
<intersection>-143 1</intersection></vsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>173,-143,173,-132.5</points>
<intersection>-143 12</intersection>
<intersection>-132.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>173,-143,211,-143</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>135.5,-132.5,173,-132.5</points>
<connection>
<GID>429</GID>
<name>IN_0</name></connection>
<intersection>173 0</intersection></hsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>223,-150.5,226.5,-150.5</points>
<connection>
<GID>435</GID>
<name>IN_0</name></connection>
<connection>
<GID>433</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>232.5,-150.5,232.5,-150.5</points>
<connection>
<GID>435</GID>
<name>OUT_0</name></connection>
<connection>
<GID>436</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>217,-144,219,-144</points>
<connection>
<GID>432</GID>
<name>N_in0</name></connection>
<connection>
<GID>430</GID>
<name>OUT</name></connection>
<intersection>217 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>217,-154,217,-144</points>
<connection>
<GID>433</GID>
<name>IN_1</name></connection>
<connection>
<GID>433</GID>
<name>IN_0</name></connection>
<intersection>-154 3</intersection>
<intersection>-144 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>217,-154,217.5,-154</points>
<connection>
<GID>434</GID>
<name>N_in3</name></connection>
<intersection>217 2</intersection></hsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-170.5,135,-170.5</points>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<connection>
<GID>439</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-171.5,142,-170.5</points>
<intersection>-171.5 1</intersection>
<intersection>-170.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-171.5,144,-171.5</points>
<connection>
<GID>440</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-170.5,142,-170.5</points>
<connection>
<GID>439</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136.5,-174.5,136.5,-173.5</points>
<intersection>-174.5 2</intersection>
<intersection>-173.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136.5,-173.5,144,-173.5</points>
<connection>
<GID>440</GID>
<name>IN_1</name></connection>
<intersection>136.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-174.5,136.5,-174.5</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<intersection>136.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133.5,-180,136,-180</points>
<connection>
<GID>442</GID>
<name>IN_0</name></connection>
<connection>
<GID>444</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>143,-181,143,-180</points>
<intersection>-181 1</intersection>
<intersection>-180 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>143,-181,144,-181</points>
<connection>
<GID>445</GID>
<name>IN_0</name></connection>
<intersection>143 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>142,-180,143,-180</points>
<connection>
<GID>444</GID>
<name>OUT_0</name></connection>
<intersection>143 0</intersection></hsegment></shape></wire>
<wire>
<ID>290</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139,-184,139,-183</points>
<intersection>-184 2</intersection>
<intersection>-183 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>139,-183,144,-183</points>
<connection>
<GID>445</GID>
<name>IN_1</name></connection>
<intersection>139 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-184,139,-184</points>
<connection>
<GID>443</GID>
<name>IN_0</name></connection>
<intersection>139 0</intersection></hsegment></shape></wire>
<wire>
<ID>291</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154.5,-185.5,154.5,-182</points>
<intersection>-185.5 9</intersection>
<intersection>-184 10</intersection>
<intersection>-182 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>150,-182,154.5,-182</points>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>152,-185.5,154.5,-185.5</points>
<connection>
<GID>446</GID>
<name>N_in0</name></connection>
<intersection>154.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>154.5,-184,159.5,-184</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<intersection>154.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>292</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-170.5,146.5,-166.5</points>
<intersection>-170.5 5</intersection>
<intersection>-166.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>146.5,-170.5,160,-170.5</points>
<connection>
<GID>448</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>133.5,-166.5,146.5,-166.5</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>293</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>150,-172.5,160,-172.5</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<intersection>152 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>152,-172.5,152,-169.5</points>
<connection>
<GID>441</GID>
<name>N_in0</name></connection>
<intersection>-172.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>294</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-178.5,167,-167</points>
<intersection>-178.5 6</intersection>
<intersection>-171.5 1</intersection>
<intersection>-169 7</intersection>
<intersection>-167 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>166,-171.5,167,-171.5</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>166,-167,167,-167</points>
<connection>
<GID>449</GID>
<name>N_in0</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>167,-178.5,176,-178.5</points>
<connection>
<GID>455</GID>
<name>IN_B_0</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>167,-169,173,-169</points>
<connection>
<GID>453</GID>
<name>IN_0</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>295</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>146.5,-188,146.5,-186</points>
<intersection>-188 6</intersection>
<intersection>-186 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>146.5,-186,159.5,-186</points>
<connection>
<GID>451</GID>
<name>IN_1</name></connection>
<intersection>146.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>133.5,-188,146.5,-188</points>
<connection>
<GID>450</GID>
<name>IN_0</name></connection>
<intersection>146.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>296</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>168.5,-187,168.5,-178.5</points>
<intersection>-187 4</intersection>
<intersection>-185 5</intersection>
<intersection>-178.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>165.5,-187,168.5,-187</points>
<intersection>165.5 7</intersection>
<intersection>168.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>165.5,-185,168.5,-185</points>
<connection>
<GID>451</GID>
<name>OUT</name></connection>
<intersection>168.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>165.5,-188,165.5,-187</points>
<connection>
<GID>452</GID>
<name>N_in0</name></connection>
<intersection>-187 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>168.5,-178.5,178,-178.5</points>
<connection>
<GID>455</GID>
<name>IN_0</name></connection>
<intersection>168.5 0</intersection>
<intersection>173 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>173,-178.5,173,-171</points>
<connection>
<GID>453</GID>
<name>IN_1</name></connection>
<intersection>-178.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>297</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-188,177,-184.5</points>
<connection>
<GID>456</GID>
<name>N_in3</name></connection>
<connection>
<GID>455</GID>
<name>OUT_0</name></connection>
<intersection>-186 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>177,-186,188.5,-186</points>
<intersection>177 0</intersection>
<intersection>188.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>188.5,-186,188.5,-183</points>
<connection>
<GID>460</GID>
<name>IN_1</name></connection>
<intersection>-186 5</intersection></vsegment></shape></wire>
<wire>
<ID>298</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196,-187,196,-175</points>
<intersection>-187 5</intersection>
<intersection>-182 6</intersection>
<intersection>-175 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>196,-175,198,-175</points>
<connection>
<GID>461</GID>
<name>IN_1</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>194.5,-187,196,-187</points>
<connection>
<GID>463</GID>
<name>N_in0</name></connection>
<intersection>196 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>194.5,-182,196,-182</points>
<connection>
<GID>460</GID>
<name>OUT</name></connection>
<intersection>196 0</intersection></hsegment></shape></wire>
<wire>
<ID>299</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>205,-177.5,205,-174</points>
<connection>
<GID>466</GID>
<name>N_in3</name></connection>
<intersection>-175 3</intersection>
<intersection>-174 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>204,-174,205,-174</points>
<connection>
<GID>461</GID>
<name>OUT</name></connection>
<intersection>205 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>205,-175,209,-175</points>
<connection>
<GID>465</GID>
<name>IN_1</name></connection>
<intersection>205 0</intersection></hsegment></shape></wire>
<wire>
<ID>300</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179.5,-170,179.5,-164.5</points>
<intersection>-170 2</intersection>
<intersection>-164.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>179.5,-164.5,188.5,-164.5</points>
<connection>
<GID>454</GID>
<name>N_in0</name></connection>
<intersection>179.5 0</intersection>
<intersection>188.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179,-170,179.5,-170</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<intersection>179.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>188.5,-166,188.5,-164.5</points>
<connection>
<GID>459</GID>
<name>IN_0</name></connection>
<intersection>-164.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>301</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>160,-180.5,160,-177.5</points>
<intersection>-180.5 10</intersection>
<intersection>-177.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>160,-180.5,188.5,-180.5</points>
<intersection>160 0</intersection>
<intersection>181 12</intersection>
<intersection>188.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>131.5,-177.5,160,-177.5</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<intersection>160 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>181,-180.5,181,-174.5</points>
<connection>
<GID>458</GID>
<name>IN_0</name></connection>
<intersection>-180.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>188.5,-181,188.5,-180.5</points>
<connection>
<GID>460</GID>
<name>IN_0</name></connection>
<intersection>-180.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>302</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>187.5,-174.5,187.5,-168</points>
<intersection>-174.5 4</intersection>
<intersection>-168 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>187.5,-168,188.5,-168</points>
<connection>
<GID>459</GID>
<name>IN_1</name></connection>
<intersection>187.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>187,-174.5,187.5,-174.5</points>
<connection>
<GID>458</GID>
<name>OUT_0</name></connection>
<intersection>187.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>303</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-173,195.5,-166</points>
<connection>
<GID>462</GID>
<name>N_in2</name></connection>
<intersection>-173 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194.5,-173,198,-173</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>194.5 3</intersection>
<intersection>195.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>194.5,-173,194.5,-167</points>
<connection>
<GID>459</GID>
<name>OUT</name></connection>
<intersection>-173 1</intersection></vsegment></shape></wire>
<wire>
<ID>304</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-173,171,-162.5</points>
<intersection>-173 12</intersection>
<intersection>-162.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>171,-173,209,-173</points>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>171 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>133.5,-162.5,171,-162.5</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>305</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,-180.5,224.5,-180.5</points>
<connection>
<GID>468</GID>
<name>OUT</name></connection>
<connection>
<GID>470</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>306</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>230.5,-180.5,230.5,-180.5</points>
<connection>
<GID>470</GID>
<name>OUT_0</name></connection>
<connection>
<GID>471</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>307</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>215,-174,217,-174</points>
<connection>
<GID>465</GID>
<name>OUT</name></connection>
<connection>
<GID>467</GID>
<name>N_in0</name></connection>
<intersection>215 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>215,-184,215,-174</points>
<connection>
<GID>468</GID>
<name>IN_1</name></connection>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<intersection>-184 3</intersection>
<intersection>-174 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>215,-184,215.5,-184</points>
<connection>
<GID>469</GID>
<name>N_in3</name></connection>
<intersection>215 2</intersection></hsegment></shape></wire>
<wire>
<ID>308</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>132.5,-202.5,134,-202.5</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<connection>
<GID>474</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>309</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141,-203.5,141,-202.5</points>
<intersection>-203.5 1</intersection>
<intersection>-202.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141,-203.5,143,-203.5</points>
<connection>
<GID>475</GID>
<name>IN_0</name></connection>
<intersection>141 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140,-202.5,141,-202.5</points>
<connection>
<GID>474</GID>
<name>OUT_0</name></connection>
<intersection>141 0</intersection></hsegment></shape></wire>
<wire>
<ID>310</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-206.5,135.5,-205.5</points>
<intersection>-206.5 2</intersection>
<intersection>-205.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-205.5,143,-205.5</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,-206.5,135.5,-206.5</points>
<connection>
<GID>472</GID>
<name>IN_0</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>311</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>132.5,-212,135,-212</points>
<connection>
<GID>477</GID>
<name>IN_0</name></connection>
<connection>
<GID>479</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>312</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-213,142,-212</points>
<intersection>-213 1</intersection>
<intersection>-212 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142,-213,143,-213</points>
<connection>
<GID>480</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>141,-212,142,-212</points>
<connection>
<GID>479</GID>
<name>OUT_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>313</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-216,138,-215</points>
<intersection>-216 2</intersection>
<intersection>-215 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-215,143,-215</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>131,-216,138,-216</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>314</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>153.5,-217.5,153.5,-214</points>
<intersection>-217.5 9</intersection>
<intersection>-216 10</intersection>
<intersection>-214 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>149,-214,153.5,-214</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<intersection>153.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>151,-217.5,153.5,-217.5</points>
<connection>
<GID>481</GID>
<name>N_in0</name></connection>
<intersection>153.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>153.5,-216,158.5,-216</points>
<connection>
<GID>486</GID>
<name>IN_0</name></connection>
<intersection>153.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>315</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-202.5,145.5,-198.5</points>
<intersection>-202.5 5</intersection>
<intersection>-198.5 6</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>145.5,-202.5,159,-202.5</points>
<connection>
<GID>483</GID>
<name>IN_0</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>132.5,-198.5,145.5,-198.5</points>
<connection>
<GID>482</GID>
<name>IN_0</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>316</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>149,-204.5,159,-204.5</points>
<connection>
<GID>475</GID>
<name>OUT</name></connection>
<connection>
<GID>483</GID>
<name>IN_1</name></connection>
<intersection>151 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>151,-204.5,151,-201.5</points>
<connection>
<GID>476</GID>
<name>N_in0</name></connection>
<intersection>-204.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>317</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>166,-210.5,166,-199</points>
<intersection>-210.5 6</intersection>
<intersection>-203.5 1</intersection>
<intersection>-201 7</intersection>
<intersection>-199 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-203.5,166,-203.5</points>
<connection>
<GID>483</GID>
<name>OUT</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>165,-199,166,-199</points>
<connection>
<GID>484</GID>
<name>N_in0</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>166,-210.5,175,-210.5</points>
<connection>
<GID>490</GID>
<name>IN_B_0</name></connection>
<intersection>166 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>166,-201,172,-201</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>166 0</intersection></hsegment></shape></wire>
<wire>
<ID>318</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145.5,-220,145.5,-218</points>
<intersection>-220 6</intersection>
<intersection>-218 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>145.5,-218,158.5,-218</points>
<connection>
<GID>486</GID>
<name>IN_1</name></connection>
<intersection>145.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>132.5,-220,145.5,-220</points>
<connection>
<GID>485</GID>
<name>IN_0</name></connection>
<intersection>145.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>319</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167.5,-219,167.5,-210.5</points>
<intersection>-219 4</intersection>
<intersection>-217 5</intersection>
<intersection>-210.5 9</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>164.5,-219,167.5,-219</points>
<intersection>164.5 7</intersection>
<intersection>167.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>164.5,-217,167.5,-217</points>
<connection>
<GID>486</GID>
<name>OUT</name></connection>
<intersection>167.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>164.5,-220,164.5,-219</points>
<connection>
<GID>487</GID>
<name>N_in0</name></connection>
<intersection>-219 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>167.5,-210.5,177,-210.5</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<intersection>167.5 0</intersection>
<intersection>172 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>172,-210.5,172,-203</points>
<connection>
<GID>488</GID>
<name>IN_1</name></connection>
<intersection>-210.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>320</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-220,176,-216.5</points>
<connection>
<GID>491</GID>
<name>N_in3</name></connection>
<connection>
<GID>490</GID>
<name>OUT_0</name></connection>
<intersection>-218 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>176,-218,187.5,-218</points>
<intersection>176 0</intersection>
<intersection>187.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>187.5,-218,187.5,-215</points>
<connection>
<GID>495</GID>
<name>IN_1</name></connection>
<intersection>-218 5</intersection></vsegment></shape></wire>
<wire>
<ID>321</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195,-219,195,-207</points>
<intersection>-219 5</intersection>
<intersection>-214 6</intersection>
<intersection>-207 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>195,-207,197,-207</points>
<connection>
<GID>496</GID>
<name>IN_1</name></connection>
<intersection>195 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>193.5,-219,195,-219</points>
<connection>
<GID>498</GID>
<name>N_in0</name></connection>
<intersection>195 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>193.5,-214,195,-214</points>
<connection>
<GID>495</GID>
<name>OUT</name></connection>
<intersection>195 0</intersection></hsegment></shape></wire>
<wire>
<ID>322</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204,-209.5,204,-206</points>
<connection>
<GID>501</GID>
<name>N_in3</name></connection>
<intersection>-207 3</intersection>
<intersection>-206 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>203,-206,204,-206</points>
<connection>
<GID>496</GID>
<name>OUT</name></connection>
<intersection>204 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>204,-207,208,-207</points>
<connection>
<GID>500</GID>
<name>IN_1</name></connection>
<intersection>204 0</intersection></hsegment></shape></wire>
<wire>
<ID>323</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>178.5,-202,178.5,-196.5</points>
<intersection>-202 2</intersection>
<intersection>-196.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>178.5,-196.5,187.5,-196.5</points>
<connection>
<GID>489</GID>
<name>N_in0</name></connection>
<intersection>178.5 0</intersection>
<intersection>187.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>178,-202,178.5,-202</points>
<connection>
<GID>488</GID>
<name>OUT</name></connection>
<intersection>178.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>187.5,-198,187.5,-196.5</points>
<connection>
<GID>494</GID>
<name>IN_0</name></connection>
<intersection>-196.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>324</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>159,-212.5,159,-209.5</points>
<intersection>-212.5 10</intersection>
<intersection>-209.5 11</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>159,-212.5,187.5,-212.5</points>
<intersection>159 0</intersection>
<intersection>180 12</intersection>
<intersection>187.5 13</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>130.5,-209.5,159,-209.5</points>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>159 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>180,-212.5,180,-206.5</points>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>-212.5 10</intersection></vsegment>
<vsegment>
<ID>13</ID>
<points>187.5,-213,187.5,-212.5</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<intersection>-212.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>325</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>186.5,-206.5,186.5,-200</points>
<intersection>-206.5 4</intersection>
<intersection>-200 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>186.5,-200,187.5,-200</points>
<connection>
<GID>494</GID>
<name>IN_1</name></connection>
<intersection>186.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>186,-206.5,186.5,-206.5</points>
<connection>
<GID>493</GID>
<name>OUT_0</name></connection>
<intersection>186.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>326</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-205,194.5,-198</points>
<connection>
<GID>497</GID>
<name>N_in2</name></connection>
<intersection>-205 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,-205,197,-205</points>
<connection>
<GID>496</GID>
<name>IN_0</name></connection>
<intersection>193.5 3</intersection>
<intersection>194.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>193.5,-205,193.5,-199</points>
<connection>
<GID>494</GID>
<name>OUT</name></connection>
<intersection>-205 1</intersection></vsegment></shape></wire>
<wire>
<ID>327</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-205,170,-194.5</points>
<intersection>-205 12</intersection>
<intersection>-194.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>170,-205,208,-205</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>132.5,-194.5,170,-194.5</points>
<connection>
<GID>499</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>328</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220,-212.5,223.5,-212.5</points>
<connection>
<GID>503</GID>
<name>OUT</name></connection>
<connection>
<GID>505</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>329</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>229.5,-212.5,229.5,-212.5</points>
<connection>
<GID>505</GID>
<name>OUT_0</name></connection>
<connection>
<GID>506</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>330</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>214,-206,216,-206</points>
<connection>
<GID>500</GID>
<name>OUT</name></connection>
<connection>
<GID>502</GID>
<name>N_in0</name></connection>
<intersection>214 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>214,-216,214,-206</points>
<connection>
<GID>503</GID>
<name>IN_1</name></connection>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<intersection>-216 3</intersection>
<intersection>-206 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>214,-216,214.5,-216</points>
<connection>
<GID>504</GID>
<name>N_in3</name></connection>
<intersection>214 2</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,890.88,1138,293.88</PageViewport></page 1>
<page 2>
<PageViewport>0,890.88,1138,293.88</PageViewport></page 2>
<page 3>
<PageViewport>0,890.88,1138,293.88</PageViewport></page 3>
<page 4>
<PageViewport>0,890.88,1138,293.88</PageViewport></page 4>
<page 5>
<PageViewport>0,890.88,1138,293.88</PageViewport></page 5>
<page 6>
<PageViewport>0,890.88,1138,293.88</PageViewport></page 6>
<page 7>
<PageViewport>0,890.88,1138,293.88</PageViewport></page 7>
<page 8>
<PageViewport>0,890.88,1138,293.88</PageViewport></page 8>
<page 9>
<PageViewport>0,890.88,1138,293.88</PageViewport></page 9></circuit>